* OPA348
*****************************************************************************
* (C) Copyright 2012 Texas Instruments Incorporated. All rights reserved.                                            
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of 
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer.
*****************************************************************************
*
* This model is subject to change without notice. Texas Instruments
* Incorporated is not responsible for updating this model.
*
*****************************************************************************
*
** Released by: Analog eLab Design Center, Texas Instruments Inc.
* Part: OPA348
* Date: 12JAN2012
* Model Type: ALL IN ONE
* Simulator: PSPICE
* Simulator Version: 16.0.0.001p
* EVM Order Number: N/A
* EVM Users Guide: N/A
* Datasheet: SBOS213D � NOVEMBER 2001 � REVISED FEBRUARY 2009
*
* Model Version: 1.0
*
*****************************************************************************
* 
* Updates:
*
* Version 1.0 : 
* Release to Web
*
*****************************************************************************
*BEGIN MODEL OPA348
*SIMULATED FEATURES:
*OPEN LOOP GAIN AND PHASE VS FREQUENCY 
*INPUT COMMON MODE REJECTION WITH FREQUENCY
*POWER SUPPLY REJECTION WITH FREQUENCY
*INPUT IMPEDANCE VS FREQUENCY 
*INPUT VOLTAGE NOISE VS FREQUENCY
*INPUT CURRENT NOISE VS FREQUENCY 
*OUTPUT VOLTAGE SWING VS OUTPUT CURRENT
*SHORT-CIRCUIT OUTPUT CURRENT
*QUIESCENT CURRENT VS SUPPLY VOLTAGE
*SLEW RATE
*SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
*LARGE SIGNAL RESPONSE
*OVERLOAD RECOVERY TIME
*INPUT BIAS CURRENT
*INPUT VOLTAGE OFFSET
*INPUT COMMON MODE RANGE
*OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS
*$
*****************************************************************************
.SUBCKT OPA348 IN+ IN- VCC VEE VOUT
V4          51 VEE 9M
V3          VCC 52 9M
IS2         54 GND_FLOAT 10P
IS1         +IN_CMRR GND_FLOAT 10P
V1          58 59 200M
V2          60 61 200M
V12         62 63 200M
V9          64 65 200M
V11         GND_FLOAT 75 10
V10         32 GND_FLOAT 10
Vor_2       78 74 800M
Vor_3       73 79 800M
EVCVS11     Vsense GND_FLOAT E GND_FLOAT  1M
EVCVS10     D GND_FLOAT C GND_FLOAT  1M
SW10        32 Over_clamp CL1 GND_FLOAT  S_VSWITCH_1
SW6         33 34 OL- GND_FLOAT  S_VSWITCH_2
SW5         35 33 GND_FLOAT OL+  S_VSWITCH_3
SW4         36 CLAW_s2 38 GND_FLOAT  S_VSWITCH_4
SW3         CLAW_s1 36 GND_FLOAT 40  S_VSWITCH_5
SW2         41 42 SC- GND_FLOAT  S_VSWITCH_6
SW1         43 41 GND_FLOAT SC+  S_VSWITCH_7
EVCVS9      46 GND_FLOAT 44 Vzo_4  1MEG
XR107       A GND_FLOAT RNOISE_FREE_0
XR107_2     46 Vzo_4 RNOISE_FREE_1
EVCVS8      B GND_FLOAT A GND_FLOAT  10U
R5          VEE VEE_A 1G 
C8          Vzo_4 GND_FLOAT 20P  
XU17        IN- P INOISE_0
XR101       0 GND_FLOAT RNOISE_FREE_2
XR102       GND_FLOAT 48 RNOISE_FREE_3
XR102_2     48 49 RNOISE_FREE_4
XR102_3     GND_FLOAT 50 RNOISE_FREE_5
XR102_4     50 PSRR RNOISE_FREE_4
XU14        GND_FLOAT Vimon VCC VEE VEE_CLP 51 VCVS_LIMIT_0
C7          GND_FLOAT AOL_p0zp1 36P 
C1          GND_FLOAT C 30P 
GVCCS10     GND_FLOAT AOL_p0zp1 D GND_FLOAT  100
XR107_3     AOL_p0zp1 GND_FLOAT RNOISE_FREE_4
XU12        VCC VEE GND_FLOAT 55 VCVS_LIMIT_1
R22         PATH+ 56 1 
R11         PATH- 57 1 
CinnCM      GND_FLOAT IN- 3P  
Cdiff       IN- IN+ 1.5P  
CinpCM      IN+ GND_FLOAT 3P  
XR107_4     CLAW_clamp GND_FLOAT RNOISE_FREE_0
XR107_5     IN+ GND_FLOAT RNOISE_FREE_6
XR107_6     GND_FLOAT IN- RNOISE_FREE_6
XR107_7     IN- IN+ RNOISE_FREE_7
XR107_8     C GND_FLOAT RNOISE_FREE_4
GVCCS2      GND_FLOAT C E GND_FLOAT  1M
XU16        Vinpins GND_FLOAT GND_FLOAT Over_clamp VCCS_LIMIT_0
C2          Over_clamp GND_FLOAT 37.5N 
XU4         VOUT Vimon GRL GND_FLOAT VCVS_GRL_0
C5          GND_FLOAT PSRR 9.43F  
C15         VCC VEE 10P  
L2          50 GND_FLOAT 1.98 
GVCCS1      GND_FLOAT PSRR VCC VEE  56.2N
CCM         49 GND_FLOAT 315F  
LCM         48 GND_FLOAT 520M  
GVCCS7      GND_FLOAT 49 +IN_CMRR GND_FLOAT  -79.4N
C4          VCC_A 0 1G 
R20         VCC VCC_A 1G 
C3          VEE_A 0 1G  
XVn11       IN+ P VNSE_0
XR104       Over_clamp GND_FLOAT RNOISE_FREE_8
XU13        +IN_CMRR P VCVS_LIMIT_2
XU11        VCC VEE 67 GND_FLOAT VCVS_LIMIT_3
XU10        VCC VEE VCC VEE VCCS_IQ_0
R32         68 PATH+ 1 
EVCVS7      61 GND_FLOAT VCC GND_FLOAT  1
XU9         68 60 IDEAL_D_0
R17         PATH+ 69 1 
XU8         59 69 IDEAL_D_0
EVCVS5      58 GND_FLOAT VEE GND_FLOAT  1
R2          70 PATH- 1 
EVCVS6      65 GND_FLOAT VCC GND_FLOAT  1
XU2         70 64 IDEAL_D_0
R3          PATH- 71 1 
XU1         63 71 IDEAL_D_0
GVCCS13     GND_FLOAT CLAW_clamp AOL_p0zp1 GND_FLOAT  10U
GVCCS14     GND_FLOAT A CLAW_clamp GND_FLOAT  10U
EVCVS2      62 GND_FLOAT VEE GND_FLOAT  1
EVCVS1      57 GND_FLOAT 54 GND_FLOAT  1
R4          VEE_CLP GND_FLOAT 100G 
R1          VCC_CLP GND_FLOAT 100G 
XU23        Vimon GND_FLOAT VCC VEE 52 VCC_CLP VCVS_LIMIT_0
C17         SC+ GND_FLOAT 1P  
C16         GND_FLOAT 38 1P  
C20         OL+ GND_FLOAT 1P
C22         GND_FLOAT CL1 1P 
R31         CL1 Over_clamp 1 
C23         GND_FLOAT Vclp 1F  
C9          72 GND_FLOAT 10P 
R30         72 Vimon 10 
C21         GND_FLOAT OL- 1P 
C19         GND_FLOAT SC- 1P 
C12         40 GND_FLOAT 1P 
R29         44 Vclp 1 
R34         Vclp 73 1K 
R33         Vclp 74 1K 
SW9         Over_clamp 75 GND_FLOAT CL1  S_VSWITCH_8
R26         42 SC- 1 
R25         43 SC+ 1 
R19         CLAW_s2 38 1 
R16         CLAW_s1 40 1 
R14         34 OL- 1 
R13         35 OL+ 1 
R12         36 CLAW_clamp 100 
R7          33 Over_clamp 10M 
R6          41 A 100 
GIsinking   VEE GND_FLOAT 76 GND_FLOAT  1M
GIsourcing  VCC GND_FLOAT 77 GND_FLOAT  1M
R23         76 GND_FLOAT 10K 
SW7         Vimon 76 72 GND_FLOAT  S_VSWITCH_9
R21         GND_FLOAT 77 10K 
SW8         Vimon 77 72 GND_FLOAT  S_VSWITCH_10
XU5         78 Vsense 35 GND_FLOAT VCVS_LIMIT_4
XU3         79 Vsense 34 GND_FLOAT VCVS_LIMIT_4
EVCVS4      56 GND_FLOAT +IN_CMRR GND_FLOAT  1
XU26        PATH+ PATH- GRL GND_FLOAT Vinpins VCCS_TG_0
XU25        PSRR GND_FLOAT 80 IN- VCVS_LIMIT_5
XU22        67 Vimon 43 GND_FLOAT VCVS_LIMIT_6
XU21        55 Vimon 42 GND_FLOAT VCVS_LIMIT_7
XU20        VEE_CLP VOUT CLAW_s2 GND_FLOAT VCVS_LIMIT_7
XU19        VCC_CLP VOUT CLAW_s1 GND_FLOAT VCVS_LIMIT_8
XR102_5     81 82 RNOISE_FREE_8
XR101_2     83 81 RNOISE_FREE_8
C6          81 0 1  
XR105       E GND_FLOAT RNOISE_FREE_8
XR103       GND_FLOAT Vinpins RNOISE_FREE_8
EVCVS34     GND_FLOAT 0 81 0  1
EVCVS29     83 0 VCC 0  1
EVCVS28     82 0 VEE 0  1
EVCVSCM     80 54 49 GND_FLOAT  1
VCCVS1_in   Vzo_4 VOUT
HCCVS1      Vimon GND_FLOAT VCCVS1_in   1K
GVCCS5      GND_FLOAT E Over_clamp GND_FLOAT  1M
EVCVS3      44 GND_FLOAT B GND_FLOAT  1

.MODEL S_VSWITCH_1 VSWITCH (RON=1 ROFF=1T VON=150 VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=1 ROFF=1T VON=1 VOFF=-1)
.MODEL S_VSWITCH_3 VSWITCH (RON=1 ROFF=1T VON=1 VOFF=-1)
.MODEL S_VSWITCH_4 VSWITCH (RON=1 ROFF=1T VON=10 VOFF=-10)
.MODEL S_VSWITCH_5 VSWITCH (RON=1 ROFF=1T VON=10 VOFF=-10)
.MODEL S_VSWITCH_6 VSWITCH (RON=1 ROFF=1T VON=10 VOFF=-10)
.MODEL S_VSWITCH_7 VSWITCH (RON=1 ROFF=1T VON=10 VOFF=-10)
.MODEL S_VSWITCH_8 VSWITCH (RON=1 ROFF=1T VON=150 VOFF=0)
.MODEL S_VSWITCH_9 VSWITCH (RON=1M ROFF=10MEG VON=-10M VOFF=0)
.MODEL S_VSWITCH_10 VSWITCH (RON=1M ROFF=10MEG VON=10M VOFF=0)
.ENDS

.SUBCKT INOISE_0 N P
XR102       87 88 RNOISE_FREE_4
GVCCS2      N P 88 0  1U
GVCCS1      0 88 89 0  565
L1          0 87 220M  
R2          89 0 1N 
.ENDS


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E5
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
*.MODEL R_RES_1 RES ( TCE=0 T_ABS=-274)
.ENDS RNOISE_FREE_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E9
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_1 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_2  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E9
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_2 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_3  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=550E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_3 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_4  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_4 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_5  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=5.63E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_5 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VC+ VC- VCC VEE VOUT+ VOUT-
.PARAM VPOS = 2
.PARAM VNEG = 0
E1 VOUT+ VOUT-  VALUE={LIMIT((V(VCC,VEE)*0.5*(0.064*V(VC+,VC-) 
+ +0.36N*V(VC+,VC-)**9)),(V(VCC,VEE)*0.5)-58M,0)}
.ENDS VCVS_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1
.PARAM VPOS = 13
.PARAM VNEG = 4.5
E1 VOUT+ VOUT- VALUE={LIMIT(5.1 + 5*(1-EXP(-1.3*(V(VC+,VC-)-2.1)))+ 
+((-2/75)*(TEMP-25)) ,VPOS,VNEG)}
.ENDS VCVS_LIMIT_1 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_6  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=20E12
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_6 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_7  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=13.33E12
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_7 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 25.12U
.PARAM IPOS = 0.01875
.PARAM INEG = -0.01875
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),IPOS,INEG)}
.ENDS VCCS_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_GRL_0  VC+ VC- VOUT+ VOUT- 
.PARAM GAIN = 1
.PARAM VPOS = 10001
.PARAM VNEG = 3000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*(3023+69.77M*((V(VC+)-V(VOUT-))/((V(VC-)-V(VOUT-))*1M))),VPOS,VNEG)}
.ENDS VCVS_GRL_0 


* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=65
* FREQ FOR 1/F VAL
.PARAM FLW=1100
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=22
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.25)/1E11} IS=1.0E-16 
* END CALC VALS
*{PWR(FLW,0.5)/1E11}
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
GR1 3 0 3 0 1N
GR2 3 0 3 0 1N
R3 3 6 1E9
GR3 3 6 3 6 1N
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
*R6 3 4 1E9
GR6 3 4 3 4 1N
R7 4 0 1E9
GR7 4 0 4 0 1N
E3 1 2 3 4 1
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE NANOV/RT-HZ


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_8  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_8 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VOUT+ VOUT-
*             
E1 VOUT+ VOUT- VALUE={1.126M+0.4U*(TEMP-25)}
.ENDS VCVS_LIMIT_2 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_3  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1
.PARAM VPOS = 13
.PARAM VNEG = 4.5
E1 VOUT+ VOUT- VALUE={LIMIT(5.1 + 5*(1-EXP(-1.3*(V(VC+,VC-)-2.1)))+ 
+((-2/75)*(TEMP-25)) ,VPOS,VNEG)}
.ENDS VCVS_LIMIT_3 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_IQ_0  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1E-6
G1 VC+ VC-  VALUE ={GAIN*(38 + 7*(1-EXP(-1.5*(V(VC+,VC-)-2.1))) + (1/10)*(TEMP-25))}
.ENDS VCCS_IQ_0 


*TG IDEAL DIODE
.SUBCKT IDEAL_D_0  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_4  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 6000
.PARAM VNEG = -6000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS VCVS_LIMIT_4 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_TG_0  VC+ VC- GRL IOUT+ IOUT-
*              
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(((V(GRL)*1u)*V(VC+,VC-)),IPOS,INEG)}
.ENDS VCCS_TG_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_5  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1
.PARAM VPOS = 20M
.PARAM VNEG = -20M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS VCVS_LIMIT_5 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_6  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1000
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS VCVS_LIMIT_6 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_7  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS VCVS_LIMIT_7 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_8  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS VCVS_LIMIT_8 