* OPA170
*****************************************************************************
* (C) Copyright 2011 Texas Instruments Incorporated. All rights reserved.                                            
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of 
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer.
*****************************************************************************
*
** Released by: Analog eLab Design Center, Texas Instruments Inc.
* Part: OPA170
* Date: 09/07/2011
* Model Type: All In One
* Simulator: TINA-TI
* Simulator Version: 9.2.30.221 SF-TI
* EVM Order Number: N/A 
* EVM Users Guide: N/A
* Datasheet: SBOS557A �AUGUST 2011�REVISED SEPTEMBER 2011
*
* Model Version: 1.0
*
*****************************************************************************
*
* Updates:
*
* Version 1.0 : Release to Web
*
*****************************************************************************
* Notes: 
*
**     Green-Lis Macromodel Architecture
*
*       OPAx170  Rev. A  by Marek Lis; 
*       August 31, 2011
*
* This macromodel has been optimized to model the AC, DC, noise, and transient response performance within 
* the device data sheet specified limits. Correct operation of this macromodel has been verified on DesignSoft
* TINA Version 9.2.30.221 SF-TI. For help with other analog simulation software, please consult the software supplier.
*
* GREEN-LIS MACRO-MODEL SIMULATED FEATURES:
*
* OPEN LOOP GAIN AND PHASE VS FREQUENCY WITH RL AND CL EFFECTS
* INPUT COMMON-MODE REJECTION VS FREQUENCY
* POWER SUPPLY REJECTION VS FREQUENCY
* INPUT IMPEDANCE VS FREQUENCY 
* OUTPUT IMPEDANCE vs OUTPUT CURRENT
* INPUT VOLTAGE NOISE VS FREQUENCY
* INPUT CURRENT NOISE VS FREQUENCY 
* OUTPUT VOLTAGE SWING FOR DIFFERENT OUTPUT CURRENTS
* SHORT-CIRCUIT OUTPUT CURRENT LIMIT
* QUIESCENT CURRENT VS SUPPLY VOLTAGE
* SETTLING TIME VS CAPACITIVE LOAD
* SLEW RATE
* SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME
* INPUT BIAS CURRENT
* INPUT BIAS OFFSET CURRENT
* INPUT VOLTAGE OFFSET
* INPUT COMMON MODE VOLTAGE RANGE
* OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS
*
* BEGIN MODEL OPA170
.SUBCKT OPA170 IN- IN+ V- V+ Vout
V7          45 8 100M
Vos         24 36 -214.1U
V11         49 50 100M
V10         51 52 100M
V6          7 57 10
V5          58 7 10
V4          54 56 800M
V1          55 53 800M
V9          69 9 2
IS2         V+ 24 8P
IS1         V+ V- 110U
IS3         41 V- -4P
V3          73 7 17
V2          7 74 20
C1          25 7 48F 
XU15        10 7 26 27 VC_RES_0
L1          28 7 800U IC=0 
R2          28 29 1 
GVCCS8      7 29 7 30  1
XR109       31 7 RNOISE_FREE_0
C3          31 7 5F
GVCCS4      7 31 21 7  1U
C2          32 7 5F 
XR109_2     32 7 RNOISE_FREE_1
GVCCS3      7 32 31 7  1M
R4          33 18 10M 
C7          34 35 3P 
C8          35 7 3P 
CinnCM      7 34 3P 
XIn11       36 34 FEMT_0
L2          37 7 200U 
XR109_3     21 7 RNOISE_FREE_0
XR109_4     38 7 RNOISE_FREE_0
XVn11       35 36 VNSE_0
XU14        39 7 40 41 VCVS_LIMIT_0
L3          42 7 200U 
R1          37 39 1 
GVCCS2      7 39 7 43  1
XU13        8 44 IDEAL_D_0
EVCVS5      45 7 V- 7  1
XR109_5     25 7 RNOISE_FREE_0
C11         38 7 48F 
XR109_6     20 7 RNOISE_FREE_1
GVCCS12     7 21 38 7  1U
XU5         10 7 V+ 11 VCVS_LIMIT_1
XU6         7 10 12 V- VCVS_LIMIT_2
C15         V+ V- 10P IC=0 
C22         7 17 1P 
R29         17 19 1 
C23         7 22 1P IC=0 
C9          46 7 10P IC=0 
R26         46 10 10 
C21         7 13 1P IC=0 
C20         7 14 1P IC=0 
C19         15 7 1P IC=0 
C17         16 7 1P IC=0 
C16         7 47 1P IC=0 
C12         48 7 1P IC=0 
R13         27 22 1 
R36         22 52 1M 
R35         22 50 1M 
SW12        53 49 15 7  S_VSWITCH_1
SW11        51 54 7 16  S_VSWITCH_2
R34         22 55 1K 
R33         22 56 1K 
SW10        58 19 17 7  S_VSWITCH_3
SW9         19 57 7 17  S_VSWITCH_4
R25         59 15 1 
R19         60 16 1 
R16         61 47 1 
R14         62 48 1 
R12         63 13 1 
R7          64 14 1 
R5          65 20 10M 
R6          66 19 10M 
R15         0 7 100MEG 
C13         20 7 5F
GVCCS1      7 20 32 7  1M
GIsinking   V- 7 67 7  1M
GIsourcing  V+ 7 68 7  1M
R23         67 7 10K 
SW7         10 67 46 7  S_VSWITCH_5
R21         7 68 10K 
SW8         10 68 46 7  S_VSWITCH_6
SW4         66 63 13 7  S_VSWITCH_7
SW3         64 66 7 14  S_VSWITCH_8
XU3         54 23 64 7 VCVS_LIMIT_3
XU1         53 23 63 7 VCVS_LIMIT_3
SW2         33 59 15 7  S_VSWITCH_9
SW1         60 33 7 16  S_VSWITCH_10
XU8         24 V+ IDEAL_D_1
XU12        V- 24 IDEAL_D_1
EVCVS6      69 7 V+ 7  1
R22         70 44 100 
EVCVS4      70 7 24 7  1
XU2         44 9 IDEAL_D_0
SW6         65 61 47 7  S_VSWITCH_11
SW5         62 65 7 48  S_VSWITCH_12
XU26        44 41 7 71 VCCS_LIMIT_0
XU4         71 7 7 19 VCCS_LIMIT_1
LPSR        72 7 800U IC=0 
XVCVSPSRR   29 7 40 34 VCVS_LIMIT_4
XU22        73 10 60 7 VCVS_LIMIT_5
XU21        74 10 59 7 VCVS_LIMIT_5
XU20        12 Vout 61 7 VCVS_LIMIT_5
XU19        11 Vout 62 7 VCVS_LIMIT_6
XU11        V- 41 IDEAL_D_1
XU10        41 V+ IDEAL_D_1
C10         18 7 5F
C5          21 7 5F 
XR109_7     18 7 RNOISE_FREE_1
GVCCS15     7 18 20 7  1M
GVCCS10     7 38 25 7  1U
R20         IN+ 35 100 
R18         IN- 34 100 
GVCCS6      7 25 23 7  1U
XR102       75 76 RNOISE_FREE_0
XR101       77 75 RNOISE_FREE_0
C6          75 0 1 IC=0 
XR105       23 7 RNOISE_FREE_0
XR104       19 7 RNOISE_FREE_2
XR103       7 71 RNOISE_FREE_0
EVCVS34     7 0 75 0  1
RPSR        72 30 1 
GVCCS11     7 30 V+ V-  1U
RCM         42 43 1 
EVCVS29     77 0 V+ 0  1
EVCVS28     76 0 V- 0  1
GVCCS7      7 43 24 7  1U
VCCVS1_in   26 Vout
HCCVS1      10 7 VCCVS1_in   1K
GVCCS5      7 23 19 7  1U
Ccc         19 7 39U
EVCVS3      27 7 18 7  1
.MODEL S_VSWITCH_1 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_4 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_5 VSWITCH (RON=1M ROFF=10MEG VON=-10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=1M ROFF=10MEG VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_8 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_9 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_10 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_11 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_12 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.ENDS


*VOLTAGE CONTROLLED RESISTOR
.SUBCKT VC_RES_0  1      2      3    4
*              VC+    VC-   RES1 RES2
ERES 3 40 VALUE = {900*(I(VSENSE) / SQRT((0.055*ABS(V(1,2))+0.055)/0.055))}
VSENSE 40 4 DC 0
.ENDS VC_RES_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * 1E6 }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * 1E3 }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_1 


* BEGIN PROG NSE FEMTO AMP/RT-HZ 
.SUBCKT FEMT_0  1 2
* BEGIN SETUP OF NOISE GEN - FEMPTOAMPS/RT-HZ
* INPUT THREE VARIABLES
* SET UP INSE 1/F
* FA/RHZ AT 1/F FREQ
.PARAM NLFF=.001
* FREQ FOR 1/F VAL
.PARAM FLWF=0.001
* SET UP INSE FB
* FA/RHZ FLATBAND
.PARAM NVRF=.001
* END USER INPUT
* START CALC VALS
.PARAM GLFF={PWR(.001,0.25)*.001/1164}
.PARAM RNVF={1.184*PWR(.001,2)}
.MODEL DVNF D KF={PWR(.001,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {PWR(.001,0.25)*.001/1164}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {1.184*PWR(.001,2)}
R5 5 0 {1.184*PWR(.001,2)}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE FEMTO AMP/RT-HZ


* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=132
* FREQ FOR 1/F VAL
.PARAM FLW=1
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=18.5
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(1,0.25)*132/1164}
.PARAM RNV={1.184*PWR(18.5,2)}
.MODEL DVN D KF={PWR(1,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {PWR(1,0.25)*132/1164}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {1.184*PWR(18.5,2)}
R5 5 0 {1.184*PWR(18.5,2)}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE NANOV/RT-HZ


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VCP VCM VOUTP VOUTM
*              
.PARAM GAIN = 1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUTP VOUTM VALUE={LIMIT(1*V(VCP,VCM),-10M,10M)}
.ENDS VCVS_LIMIT_0 


*TG IDEAL DIODE
.SUBCKT IDEAL_D_0  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VCP VCM VOUTP VOUTM
*              

E1 VOUTP VOUTM TABLE {ABS(V(VCP,VCM))} = (0, 0.01) (5, 0.5) (8.5, 1.0) (16.9, 2.5)
.ENDS VCVS_LIMIT_1 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VCP VCM VOUTP VOUTM
*              

E1 VOUTP VOUTM TABLE {ABS(V(VCP,VCM))} = (0, 0.01) (5, 0.25) (8, 0.5) (19.9, 1.5) 
.ENDS VCVS_LIMIT_2 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_3  VCP VCM VOUTP VOUTM
*              
.PARAM GAIN = 100
.PARAM VPOS = 6000
.PARAM VNEG = -6000
E1 VOUTP VOUTM VALUE={LIMIT(100*V(VCP,VCM),-6000,6000)}
.ENDS VCVS_LIMIT_3 


*TG IDEAL DIODE
.SUBCKT IDEAL_D_1  A C
D1 A C DNOM 
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_1 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VCP VCM IOUTP IOUTM
*              
.PARAM GAIN = 100U
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUTP IOUTM VALUE={LIMIT(100U*V(VCP,VCM),-.5,.5)}
.ENDS VCCS_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_1  VCP VCM IOUTP IOUTM
*              
.PARAM GAIN = 3.2
.PARAM IPOS = 15.6
.PARAM INEG = -15.6
G1 IOUTP IOUTM VALUE={LIMIT(3.2*V(VCP,VCM),-15.6,15.6)}
.ENDS VCCS_LIMIT_1 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_4  VCP VCM VOUTP VOUTM
*              
.PARAM GAIN = -1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUTP VOUTM VALUE={LIMIT(-1*V(VCP,VCM),-10M,10M)}
.ENDS VCVS_LIMIT_4 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_5  VCP VCM VOUTP VOUTM
*              
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUTP VOUTM VALUE={LIMIT(100*V(VCP,VCM),-5000,5000)}
.ENDS VCVS_LIMIT_5 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_6  VCP VCM VOUTP VOUTM
*             
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUTP VOUTM VALUE={LIMIT(100*V(VCP,VCM),-5000,5000)}
.ENDS VCVS_LIMIT_6 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_2  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E4
ERES 1 3 VALUE = { I(VSENSE) * 1E4 }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_2 


.END
