*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG
*SIMULATOR=PSPICE
*DATE=25/02/2009
*VERSION=1
*PIN_ORDER         D G S
*
.SUBCKT ZXMP6A17E6 1 2 3
M11 20 21 22 22 Ppmod1 L=1.4E-6 W=1.25
M12 22 21 22 20 Npmod1 L=1.4E-6 W=0.95
RG1 21 27 2.8
RIN1 21 22 1E9
RD1 20 24 Rpmod1 0.028
RS1 22 23 Rpmod1 0.068
RL1 23 24 7E9
C1 21 22 160E-12
D1 24 23  Dpmod1
LD1 1 24 0.3E-9
LG1 2 27 1.2E-9
LS1 3 23 1.2E-9
.MODEL Ppmod1 PMOS (LEVEL=3 TOX=8.6E-8 NSUB=8E15
+VTO=-2.18 KP=3.5E-5 NFS=3.5E11 KAPPA=0.016 IS=1E-15 N=10)
.MODEL Npmod1 NMOS (LEVEL=3 TOX=8.6E-8 NSUB=6.5E15 
+TPG=-1 IS=1E-15 N=10)
.MODEL Dpmod1 D (IS=2E-12 RS=0.02 IKF=0.1 TRS1=1.5e-3 CJO=85e-12 
+M=0.43 VJ=0.41 TT=3.2e-8  BV=66)
.MODEL Rpmod1 RES (TC1=4.6e-3 TC2=8E-6)
.ENDS
*
*$