**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: FQT7N10
** 100V N-Channel MOSFET and TO-223
** Model Type: BSIM3V3
**-------------------------------------------------------------------------------
.SUBCKT FQT7N10 2 1 3
*Nom Temp=25 deg C
Dbody 7 5    DbodyMOD
Dbreak 5 11  DbreakMOD
Ebreak 11 7 17 7 110
Lgate 1 9    1.566e-9
Ldrain 2 5   1.44e-9
Lsource 3 7  1.874e-9
RLgate 1 9   15.7
RLdrain 2 5  14.4
RLsource 3 7 18.7
Rgate 9 6    1.5
It 7 17      1
Rbreak 17 7  RbreakMOD 1
.MODEL RbreakMOD RES (TC1=1.01e-3 TC2=-1.14e-6)
.MODEL DbodyMOD D (IS=2.85e-13 N=1      RS=3.62e-2  TRS1=3.8e-3 TRS2=1.0e-6
+ CJO=2.84e-10     M=0.24      VJ=0.45  TT=6.25e-8  XTI=3       EG=1.32)
.MODEL DbreakMOD D (RS=100e-3 TRS1=1.0e-3 TRS2=1e-6)
Rdrain 5 16 RdrainMOD 0.22
.MODEL RdrainMOD RES (TC1=7.2e-3 TC2=2.16e-5)
M_BSIM3 16 6 7 7 Bsim3 W=0.25 L=2.0e-6 NRS=1
.MODEL  Bsim3 NMOS (LEVEL=7 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=780e-10     XJ=1.4e-6      NCH=1.3e17      UA=8.8e-9
+ U0=700          VSAT=1.0e5     DROUT=1.0
+ DELTA=0.1       PSCBE2=0       RSH=1.09e-3
+ VTH0=2.83       VOFF=-0.1      NFACTOR=1.1
+ LINT=5.4e-7     DLC=5.4e-7     
+ CGSO=4.5e-10    CGSL=0         CGDO=9.65e-13
+ CGDL=1.08e-9    CJ=0           CF=0
+ CKAPPA=0.2      KT1=-1.32      KT2=0
+ UA1=6.0e-10     NJ=10
.ENDS
