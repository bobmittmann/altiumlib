.SUBCKT BSP250 1 2 3
* 1=drain  2=gate  3=source
Cgs  6 3 216e-12
Cgd1 6 4 529e-12
Cgd2 1 4 50e-12
M1 5 6 3 3 MOST1
M2 4 6 5 3 MOST2
D1 1 3 Dbody
Rd 5 1 Rtemp 25e-3
Rg 2 6 50
.MODEL MOST1 PMOS(Level=3 Vto=-1.6 Kp=9.5e-8 Eta=1e-5 W=1 L=0.1e-6
+                Rs=0 Rd=0 Ld=0 Wd=0 Uo=500 Vmax=4e7
+                Xj=5e-7 Kappa=0.08 Nfs=3e12 Theta=5e-3 Tpg=1
+                Cgbo=0 Cgso=0 Cgdo=0 Delta=0.1 Is=0)
.MODEL MOST2 PMOS(Level=3 Vto=3.8 Kp=9.5e-8 Eta=1e-5 W=1.5e-4 L=0.1e-6
+                Rs=0 Rd=0 Ld=0 Wd=0 Uo=500 Vmax=0
+                Xj=0 Kappa=0.2 Nfs=0 Theta=0 Tpg=1
+                Cgbo=0 Cgso=0 Cgdo=0 Delta=0 Is=0)
.MODEL Dbody D(Is=1e-14 N=1 Rs=190e-3 Ikf=1e3 Cjo=0 M=0.5 Vj=0.4
+                Bv=30 Ibv=10e-6 Tt=230e-9)
.MODEL Rtemp RES(TC1=4.15e-3 TC2=2e-6)
.ENDS
