.SUBCKT SMT1N  2  3  50  60
* SCHMITT-TRIGGER INPUT FOR LV14 CMOS INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MLVPEN W=20U L=2.0U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MLVNEN W=35U L=2.0U AD=140P AS=140P PD=50U PS=35U
MP2 5  4 50 50  MLVPEN W=36U L=2.0U AD=140P AS=140P PD=50U PS=35U
MN2 6  4 60 60  MLVNEN W=16U L=2.0U AD= 70P AS= 70P PD=15U PS=17U
MP3 3  4  5 50  MLVPEN W=44U L=4.0U AD=220P AS=220P PD=60U PS=44U
MN3 3  4  6  6  MLVNEN W=17U L=2.0U AD= 70P AS= 70P PD=15U PS=16U
MP4 5  3 60 50  MLVPEN W=36U L=2.0U AD=150P AS=150P PD=60U PS=36U
MN4 6  3 50  6  MLVNEN W= 6U L=4.0U AD= 25P AS= 25P PD=10U PS= 6U
.MODEL MLVNEN NMOS LEVEL=3 KP=65.0E-6 VTO=0.46 TOX=30.0E-9 NSUB=2.8E15 GAMMA=0.94 PHI=0.65 VMAX=150E3 RS=30 RD=30 XJ=0.11E-6 LD=0.4E-6 DELTA=0.315 THETA=0.054 ETA=0.015 KAPPA=0.0
.MODEL MLVPEN PMOS LEVEL=3 KP=20.3E-6 VTO=-0.61 TOX=30.0E-9 NSUB=3.3E16 GAMMA=0.92 PHI=0.65 VMAX=970E3 RS=60 RD=60 XJ=0.63E-6 LD=0.15E-6 DELTA=2.24 THETA=0.108 ETA=0.322 KAPPA=0.0
.ENDS

.SUBCKT INVN   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MLVPEN W=364U L=2.0U AD=500P  AS=500P PD=10U PS=430U
MN1 3  2 60 60  MLVNEN W=184U L=2.0U AD=275P  AS=275P PD=10U PS=270U
.MODEL MLVNEN NMOS LEVEL=3 KP=65.0E-6 VTO=0.46 TOX=30.0E-9 NSUB=2.8E15 GAMMA=0.94 PHI=0.65 VMAX=150E3 RS=30 RD=30 XJ=0.11E-6 LD=0.4E-6 DELTA=0.315 THETA=0.054 ETA=0.015 KAPPA=0.0
.MODEL MLVPEN PMOS LEVEL=3 KP=20.3E-6 VTO=-0.61 TOX=30.0E-9 NSUB=3.3E16 GAMMA=0.92 PHI=0.65 VMAX=970E3 RS=60 RD=60 XJ=0.63E-6 LD=0.15E-6 DELTA=2.24 THETA=0.108 ETA=0.322 KAPPA=0.0
.ENDS

.SUBCKT OUTPN 2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MLVPEN W=360U L=2.0U AD=400P AS=400P PD=10U PS=180U
MN1 3 4 60 60  MLVNEN W=140U L=2.0U AD=200P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MLVPEN W=360U L=2.0U AD=400P AS=400P PD=10U PS=180U
MN2 3 5 60 60  MLVNEN W=140U L=2.0U AD=200P AS=200P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MLVPEN W=360U L=2.0U AD=400P AS=400P PD=10U PS=180U
MN3 3 6 60 60  MLVNEN W=140U L=2.0U AD=200P AS=200P PD=10U PS=130U
.MODEL MLVNEN NMOS LEVEL=3 KP=65.0E-6 VTO=0.46 TOX=30.0E-9 NSUB=2.8E15 GAMMA=0.94 PHI=0.65 VMAX=150E3 RS=30 RD=30 XJ=0.11E-6 LD=0.4E-6 DELTA=0.315 THETA=0.054 ETA=0.015 KAPPA=0.0
.MODEL MLVPEN PMOS LEVEL=3 KP=20.3E-6 VTO=-0.61 TOX=30.0E-9 NSUB=3.3E16 GAMMA=0.92 PHI=0.65 VMAX=970E3 RS=60 RD=60 XJ=0.63E-6 LD=0.15E-6 DELTA=2.24 THETA=0.108 ETA=0.322 KAPPA=0.0
.ENDS

.SUBCKT INVSMT  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    SMT1N
XINV  25  30  50  60    INVN
XOUTP 30  40  50  60    OUTPN
L1  80  50   3.54NH
L2  60  90   3.54NH
L3   2  20   3.54NH
L4  40   3   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


