*SRC=DMP3020LSS;DI_DMP3020LSS;MOSFETs P;Enh;30.0V 12.0A 25.0mohms  Diodes Inc MOSFET
*SYM=POWMOSP
.SUBCKT DI_DMP3020LSS   10 20 30
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  10.9m
RS  40  3  1.62m
RG  20  2  76.7
CGS  2  3  179p
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  347p
R1  13  0  1.00
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1.00
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.50n
.MODEL DMOS PMOS(LEVEL=3 VMAX=62.5k THETA=80.0m
+ ETA=450u VTO=-2.00 KP=23.3
.MODEL DCGD D (CJO=347p VJ=0.600 M=0.680
.MODEL DSUB D (IS=49.8n N=1.50 RS=29.2m BV=30.0
+ CJO=92.5p VJ=0.800 M=0.420 TT=196n
.MODEL DLIM D (IS=100U)
.ENDS

