* ------------------------------
* Connections
*      1  = Y1  (NO)
*      2  = GND
*      3  = Y0  (NC)
*      4  = Z
*      5  = VCC
*      6  = S
*****************

.SUBCKT 74LVC1G3157 1 2 3 4 5 6
X1 1 3 4 6 5 2 ANALOG_SW_SPDT
.ENDS


*****************
* Connections
*      1  = NO
*      2  = NC
*      3  = CO (Common)
*      4  = SEL
*      5  = VCC
*      6  = GND
*****************

.SUBCKT ANALOG_SW_SPDT 1 2 3 4 5 6
S1 1 3 4 6 SMOD1
S2 2 3 4 6 SMOD2
*SUPPLY CURRENT
RSUPP 5 3 90MEG
*ANALOG SIGNAL RANGES
DCOM1 3 5 DX
DCOM2 6 3 DX
DNO1 1 5 DX
DNO2 6 1 DX
DNC1 2 5 DX
DNC2 6 2 DX
*CHARGE-INJECTION
CNOIN 4 1  10P
CNCIN 4 2  10P
CCOMIN 4 3 10P
*FREQUENCY RESPONSE OF OFF-ISOLATION
CNOI 1 3 5.65P
CNCI 2 3 5.65P
*MODELS USED
.MODEL SMOD1 VSWITCH(RON=6.5 ROFF=62.946E6 VON=1.4 VOFF=0.5)
.MODEL SMOD2 VSWITCH(RON=6.5 ROFF=62.946E6 VON=0.5 VOFF=1.4)
.MODEL DX D(IS=1E-18 N=0.001)
.ENDS
*****************

