*SRC=DMN3115UDM;DI_DMN3115UDM;MOSFETs N;Enh;30.0V 3.20A 60.0mohms  Diodes Inc MOSFET
.SUBCKT DI_DMN3115UDM   10 20 30
*     TERMINALS:  D  G  S
M1   10  20  30  30  DMOS L=1U W=1U
.MODEL DMOS NMOS( LEVEL=1 VTO=1.00 KP=10.7  GAMMA=1.24
+ PHI=.75  LAMBDA=50.9u RD=8.40m RS=8.40m
+ IS=1.60p  PB=0.800 MJ=0.460 CBD=76.2p
+ CBS=91.4p  CGSO=648n CGDO=540n CGBO=3.57u  )
.ENDS
*   -- Assumes default L=100U W=100U --

