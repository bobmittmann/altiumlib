* BEGIN MODEL LMV651
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THRU
* THE SUPPLY RAILS, OUTPUT SWING VS IO, OUTPUT CURRENT LIMIT,
* OPEN LOOP GAIN AND PHASE, SLEW RATE, COMMON MODE REJECTION
* WITH FREQ EFFECTS, POWER SUPPLY REJECTION WITH FREQ EFFECTS,
* INPUT VOLTAGE NOISE WITH 1/F, INPUT CURRENT NOISE, INPUT
* CAPACITANCE, INPUT BIAS CURRENT, INPUT COMMON MODE RANGE,
* INPUT OFFSET, HIGH CLOAD EFFECTS, AND QUIESCENT CURRENT
* VS VOLTAGE AND TEMPERATURE.
*///////////////////////////////////////////////////////////////
* MODEL TEMP RANGE IS -40 TO +125 DEG C. 
* NOTE THAT MODEL IS FUNCTIONAL OVER THIS	RANGE BUT NOT ALL
* PARAMETERS TRACK THOSE OF THE REAL PART.
*////////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  1   3   5  2  4
.SUBCKT LMV651 1 3 5 2 4
Q12 6 7 8 QP
Q13 9 9 10 QP
Q14 11 11 9 QP
Q15 8 12 10 QP
Q17 13 8 14 QOP
Q18 15 15 16 QN
Q19 16 16 17 QN
Q20 6 18 19 QN
Q21 20 6 21 QON
Q22 8 15 6 QN
R10 18 22 100
R11 12 23 100
R12 14 5 50
R13 2 21 4
G1 6 19 24 25 -2E-4
R16 24 26 100
C2 26 4 17E-12
R17 7 11 50
R18 19 17 4
D5 4 5 DD
D6 2 4 DD
E2 19 0 2 0 1
E3 10 0 5 0 1
I12 5 2 105E-6
G4 24 25 27 28 2E-3
R40 24 25 9E5
E14 25 19 10 19 0.5
D11 24 10 DD
D12 19 24 DD
R41 20 4 2
R42 4 13 4
Q23 8 29 10 QP
Q24 15 30 10 QP
Q25 6 31 19 QN
Q26 7 32 19 QN
Q33 33 34 10 QP
R45 35 36 1
R46 37 36 1
R47 38 39 7E3
R49 19 27 425
R50 19 28 425
R51 40 41 7E3
Q35 41 41 42 QP
Q37 42 42 41 QN
D13 42 10 DD
D14 41 10 DD
D15 43 42 DD
D16 43 41 DD
V10 39 42 -0.07E-3
D17 44 0 DIN
D18 45 0 DIN
I14 0 44 0.1E-3
I15 0 45 0.1E-3
C13 38 0 3E-12
C14 3 0 3E-12
D19 46 0 DVN
D20 47 0 DVN
I16 0 46 0.1E-3
I17 0 47 0.1E-3
E15 40 3 46 47 1.75
G5 38 40 44 45 3.6E-5
E16 49 0 10 0 1
E17 50 0 19 0 1
E18 51 0 52 0 1
R56 49 53 1E6
R57 50 54 1E6
R58 51 55 1E6
R59 0 53 100
R60 0 54 100
R61 0 55 100
E19 56 1 55 0 -47E-3
R62 57 52 1E3
R63 52 58 1E3
C15 49 53 1E-12
C16 50 54 1E-12
C17 51 55 70E-12
E20 59 56 54 0 0.25
E21 38 59 53 0 -0.20
C19 27 28 8E-12
G6 34 10 60 0 0.68E-6
G7 29 10 60 0 3.4E-7
G8 30 10 60 0 1.45E-7
G9 19 31 60 0 1.7E-7
G10 19 32 60 0 7.25E-8
R64 0 60 1E12
R132 4 24 1E8
I18 38 0 80E-9
I19 3 0 80E-9
V53 43 19 0.07
V54 33 36 0.1
G12 38 40 61 0 8E-6
R136 0 61 12E3
R137 0 61 12E3
R138 1 56 1E9
R139 56 59 1E9
R140 59 38 1E9
E54 58 0 38 0 1
E55 57 0 40 0 1
C23 38 40 0.25E-12
E72 22 19 21 2 3.5
E73 23 10 14 10 0.75
M61 28 42 35 35 MIP L=2U W=150U
M62 27 41 37 37 MIP L=2U W=150U
V55 60 0 1
R141 2 5 1E6
G13 5 2 62 0 -2E-4
I20 0 63 1E-3
D21 63 0 DD
V56 63 62 0.65
R143 0 62 1E6
.MODEL QON NPN VAF=40
.MODEL QOP PNP VAF=40
.MODEL MIP PMOS KP=600U VTO=-0.7
.MODEL DD D
.MODEL QN NPN
.MODEL QP PNP
.MODEL DVN D KF=0.7E-16
.MODEL DIN D KF=8E-17
.ENDS
* END MODEL LMV651
