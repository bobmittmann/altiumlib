*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG
*SIMULATOR=PSPICE
*DATE=25/02/09
*VERSION=1
*PIN_ORDER         D G S
*
.SUBCKT ZXMN10A08G 1 2 3
M11 20 21 22 22 Nnmod1 L=1E-6 W=0.6
M12 22 21 22 20 Pnmod1 L=1.5E-6 W=0.45
RG1 21 27 3.2
RIN1 21 22 1E12
RD1 20 24 Rnmod1 0.14
RS1 22 23 1E-6
RL1 23 24 10E9
C11 21 22 65E-12
C12 20 21 10E-12
D1 23 24  Dnmod1
LD1 1 24 1.0E-9
LG1 2 27 2.3E-9
LS1 3 23 2.3E-9
.MODEL Nnmod1 NMOS (LEVEL=3 TOX=5E-8 NSUB=2E17 VTO=4.05
+KP=18E-5 RS=.07 NFS=2E12 KAPPA=0.06 UO=650 IS=1E-15 N=10)
.MODEL Pnmod1 PMOS (LEVEL=3 TOX=15E-8 NSUB=2E15
+TPG=-1 IS=1E-15 N=10)
.MODEL Dnmod1 D (IS=2E-12 RS=.02 IKF=0.06 TRS1=1.5e-3
+CJO=120e-12 BV=110)
.MODEL Rnmod1 RES (TC1=9.5e-3 TC2=2.5E-5)
.ENDS ZXMN10A08G
*
*$