* BEGIN MODEL LMV641
* Rev. A October-2007
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
*MODEL KEY FEATURES INCLUDE:
* OUTPUT SWING, OPEN LOOP GAIN AND PHASE, SLEW RATE, 
* COMMON MODE REJECTION vs FREQUENCY, POWER SUPPLY REJECTION vs FREQUENCY,
* INPUT VOLTAGE NOISE WITH 1/F, OUTPUT SATURATION VOLTAGE,
* INPUT CAPACITANCE, INPUT BIAS CURRENT, INPUT COMMON MODE RANGE, 
* INPUT OFFSET VOLTAGE, QUIESCENT SUPPLY CURRENT.
*//////////////////////////////////////////////////////////////////////
*MODEL TEMP RANGE IS +25 DEG C (ROOM TEMP ONLY).
* Vsupply = +/-5V
* DEVICE PINOUT ORDER  +IN -IN +V -V OUT
* DEVICE PIN NUMBER     1   3   5  2  4 
*//////////////////////////////////////////////////////////////////
* Node Assignments
*              noninverting input
*              | inverting input
*              | | positive supply
*              | | |  negative supply
*              | | |  |  output
*              | | |  |  |
*              | | |  |  |
.SUBCKT LMV641 1 2 99 50 45
*
*  INPUT STAGE
*
Q1    5  7  3 PIX
Q2    6  2  4 PIX
RC1   5 50 4E3
RC2   6 50 4E3
RE1   3 10 68.5
RE2   4 10 68.5
I1   99 10 100E-6
C1    5  6 8.44E-13
D1    3  8 DX
V1   99  8  1.5
EOS   7  1 POLY(5) (73,98) (22,98) (81,98) (80,98) (83,98) 0.4E-3 1 1 1 1 1
IOS   1  2 1.1E-9

*
*CMRR Network
*
E1  72 98 POLY(2) (1,98) (2,98) 0 5E-01 5E-01
R10 72 73 1.59E+02
R20 73 98 1.59E-03
C10 72 73 1.00E-06
*
* PSRR Network
*
EPSY 21 98 POLY(1) (99,50) -1.2E-02 1
RPS1 21 22 1.59E+2
RPS2 22 98 1.59E-3
CPS1 21 22 1.00E-06

* VOLTAGE NOISE REFERENCE OF 15nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 14
RN2 81 98 1
*
* FLICKER NOISE CORNER 
*
DFN 82 98 DNOISE
VFN 82 98 DC 0.6551
HFN 83 98 POLY(1) VFN 1.00E-03 1.00E+00
RFN 83 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) -7.65E-03 3E-05
EVP  97 98 (99,50) 0.5
EVN  51 98 (50,99) 0.5
*

*
* GAIN STAGE
*
G1   98 30 POLY(1) (5,6)  0 17E-3
R1   30 98 1E6
CF   30 31 1.7E-9
Rz   31 45 2
D5   30 97 DX
D6   51 30 DX
*
* RAIL-TO-RAIL OUTPUT STAGE
*
Q5   45 41 99 POUT
Q6   45 43 50 NOUT
EB1  99 40 POLY(1) (98,30) 0.7745 1
EB2  42 50 POLY(1) (30,98) 0.7745 1
RB1  40 41 2.4e2
RB2  42 43 2.4e2
D7   46 99 DX
D8   47 43 DX
V5   46 41 0.5
V6   47 50 0.5
*

.MODEL PIX PNP (BF=625,IS=1E-16,VAF=130)
.MODEL POUT PNP (BF=625,IS=1E-15,VAF=200)
.MODEL NOUT NPN (BF=100,IS=1E-15,VAF=200)
.MODEL DX D(IS=1E-16,RS=5)
.MODEL DNOISE D(IS=1E-14,KF=2.25E-13)
.ENDS 
* END MODEL LMV641

