*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG
*SIMULATOR=PSPICE
*DATE=25/02/2009
*VERSION=3
*PIN_ORDER         D G S
*
.SUBCKT ZXMP3A16G 1 2 3
M11 20 21 22 22 Ppmod1 L=1.2E-6 W=1.67
M12 22 21 22 20 Npmod1 L=1.4E-6 W=1.4
RG1 21 27 2.0
RIN1 21 22 1E10
RD1 20 24 Rpmod1 0.0085
RS1 22 23 Rpmod1 0.025
RL1 23 24 3E9
C11 21 22 600E-12
C12 20 21 25E-12
D1 24 23  Dpmod1
LD1 1 25 1.0E-9
LG1 2 27 2.3E-9
LS1 3 23 2.3E-9
.MODEL Ppmod1 PMOS (LEVEL=3 TOX=7.5E-8 NSUB=1.5E16 VTO=-1.87
+KP=1.35E-5 NFS=4.5E11 KAPPA=0.06 IS=1E-15 N=10)
.MODEL Npmod1 NMOS (LEVEL=3 TOX=7.5E-8 NSUB=2E16
+TPG=-1 IS=1E-15 N=10)
.MODEL Dpmod1 D (IS=2.4E-12 RS=.016 IKF=0.2 TRS1=1.5e-3
+CJO=590e-12  BV=33 TT=16e-9)
.MODEL Rpmod1 RES (TC1=3.13e-3 TC2=4E-6)
.ENDS
*
*$
