*
*Zetex ZXMN2B03E6 Spice Model v1.0 Last Revised 7/12/07
*
.SUBCKT ZXMN2B03E6 30 40 50
*------connections-------D-G-S
M1 6 2 5 5 Nmod L=1.16E-6 W=1.83
M2 5 2 5 6 Pmod L=1.2E-6 W=0.67
RG 4 22 1.5
RIN 2 5 1E12
RD 3 6 Rmod1 0.015
RL 3 5 3E9
C1 2 5 10E-12
C2 3 4 3E-12
D1 5 3  Dmod1
Rt 5 61 Rmod2 1
Vt 61 62 1
It 5 62 1
Et 2 22  62 5 1
LD 3 30 0.5E-9
LG 4 40 1.0E-9
LS 5 50 1.0E-9
.MODEL Nmod NMOS (LEVEL=3 TOX=3.5E-8 NSUB=1E17 VTO=0.8
+KP=7E-5 RS=.020 NFS=1E11 KAPPA=0.06 IS=1E-15 N=10)
.MODEL Pmod PMOS (LEVEL=3 TOX=3.5E-8 NSUB=4.1E16
+TPG=-1 IS=1E-15 N=10)
.MODEL Dmod1 D (IS=1E-11 RS=.05 IKF=.5 TT=0.6E-8
+CJO=200e-12  BV=23)
.MODEL Rmod1 RES (TC1=8e-3 TC2=0.9E-5)
.MODEL Rmod2 RES (TC1=-1.2e-3 TC2=-1E-6)
.ENDS ZXMN2B03E6
*
*$
*
*                (c)  2007 Zetex Semiconductors plc
*
*   The copyright in these models  and  the designs embodied belong
*   to Zetex Semiconductors plc (" Zetex ").  They  are  supplied
*   free of charge by Zetex for the purpose of research and design
*   and may be used or copied intact  (including this notice)  for
*   that purpose only.  All other rights are reserved. The models
*   are believed accurate but  no condition  or warranty  as to their
*   merchantability or fitness for purpose is given and no liability
*   in respect of any use is accepted by Zetex, its distributors
*   or agents.
*
*   Zetex Semiconductors plc, Zetex Technology Park, Chadderton,
*   Oldham, United Kingdom, OL9 9LL

