*---------- DMG2307L Spice Model ----------
.SUBCKT DMG2307L 10 20 30
*     TERMINALS:  D  G  S
M1 1 2 3 3  PMOS  L = 1E-006  W = 1E-006
RD 10 1 0.04307
RS 30 3 0.001
RG 20 2 17.1
CGS 2 3 3.339E-010
EGD 12 30 2 1 1
VFB 14 30 0
FFB 2 1  VFB 1
CGD 13 14 3.9E-010
R1 13 30 1
D1 13 12  DLIM
DDG 14 15  DCGD
R2 12 15 1
D2 30 15  DLIM
DSD 10 3  DSUB
.MODEL PMOS PMOS  LEVEL = 3  U0 = 400  VMAX = 1E+006  ETA = 0.001
+ TOX = 6E-008  NSUB = 1E+016  KP = 8.459  KAPPA = 9.123  VTO = -1.527
.MODEL DCGD D  CJO = 1.701E-010  VJ = 0.4656  M = 0.372
.MODEL DSUB D  IS = 5E-010  N = 1.421  RS = 0.05533  BV = 33  CJO = 2.821E-011  VJ = 0.5166  M = 0.4868
.MODEL DLIM D  IS = 0.0001
.ENDS
*Diodes DMG2307L Spice Model v1.0 Last Revised 2011/10/28
