*
*NZH12B
*
*NXP Semiconductors
*
*Single Zener diode
*
*
*
*
*
*
*IR    = 0,04�A @ VR = 9V
*
*Vzmax = 12,03V @ IZ = 10mA
*
*
*
*
*
*
*
*Package pinning does not match Spice model pinning.
*Package: SOD123F
*
*Package Pin 1: Cathode
*Package Pin 2: Anode
*
*
*
*
*Simulator: SPICE3
*
*******************************************
*#
.SUBCKT NZH12B 1 2
*
*The resistor R1 and the diode D2 do not reflect
*physical devices but improve
*only modeling in the reverse
*mode of operation.
*
R1 1 2 1E+012
D1 1 2 DIODE1
D2 1 2 DIODE2
*
.MODEL DIODE1 D
+ IS = 1.5E-015
+ N = 2
+ BV = 11.72
+ IBV = 0.01
+ RS = 0.324
+ CJO = 4.25E-011
+ VJ = 0.51
+ M = 0.31
+ FC = 0.5
+ TT = 0
+ EG = 1.1
+ XTI = 3
.MODEL DIODE2 D
+ IS = 2E-016
+ N = 1
+ RS = 0.4
.ENDS
*
