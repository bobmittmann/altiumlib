* TLV271
*****************************************************************************
* (C) Copyright 2011 Texas Instruments Incorporated. All rights reserved.                                            
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of 
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer.
*****************************************************************************
*
* This model is subject to change without notice. Texas Instruments
* Incorporated is not responsible for updating this model.
*
*****************************************************************************
*
** Released by: Analog eLab Design Center, Texas Instruments Inc.
* Part: TLV271
* Date: 13JUN2011
* Model Type: ALL IN ONE
* Simulator: PSPICE
* Simulator Version: 16.0.0.p001
* EVM Order Number: N/A
* EVM Users Guide: N/A
* Datasheet: SLOS351D - MARCH 2001 - REVISED FEBRUARY 2004
*
* Model Version: 1.0
*
*****************************************************************************
* 
* Updates:
*
* Version 1.0 : 
* Release to Web
*
*****************************************************************************
*
*     connections:         non-inverting input
*                          |  inverting input
*                          |  |  positive power supply
*                          |  |  |  negative power supply
*                          |  |  |  |   output
*                          |  |  |  |   |
.subckt amp_tlv27x_highVdd 1 2 3 4 5
*
c1 11 12 457.48E-15
c2 6 7 5.0000E-12
css 10 99 1.1431E-12
dc 5 53 dy
de 54 5 dy
dlp 90 91 dx
dln 92 90 dx
dp 4 3 dx
egnd 99 0 poly(2) (3,0) (4,0) 0 .5 .5
fb 7 99 poly(5) vb vc ve vlp vln 0 176.02E6 -1E3 1E3 180E6 -180E6
ga 6 0 11 12 16.272E-6
gcm 0 6 10 99 6.8698E-9
iss 10 4 dc 1.3371E-6
hlim 90 0 vlim 1K
j1 11 2 10 jx1
J2 12 1 10 jx2
r2 6 9 100.00E3
rd1 3 11 61.456E3
rd2 3 12 61.456E3
ro1 8 5 10
ro2 7 99 10
rp 3 4 150.51E3
rss 10 99 149.58E6
vb 9 0 dc 0
vc 3 53 dc .78905
ve 54 4 dc .78905
vlim 7 8 dc 0
vlp 91 0 dc 14.200
vln 0 92 dc 14.200
.model dx D(Is=800.00E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx1 NJF(Is=500.00E-15 Beta=198.03E-6 Vto=-1)
.model jx2 NJF(Is=500.00E-15 Beta=198.03E-6 Vto=-1)
.ends
*END TLV272
