.SUBCKT MCP6471 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6471
*
* Revision History:
*      REV A: 01-Dec-12, Created model      
*
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Vos distribution, Ib distribution for Monte Carlo
*      Distortion (detailed non-linear behavior)
*      Some Temperature analysis
*      Process variation
*      Behavior outside normal operating region    
*
* Input Stage
V10  3 10 -210M
R10 10 11 69.0K
R11 10 12 69.0K
G10 10 11 10 11 1.44M
G11 10 12 10 12 1.44M
C11 11 12 115E-15
C12  1  0 6.00P
E12 71 14 VALUE { 65.0U + V(20) * 3.94 + V(21) * 3.94 + V(22) * 3.94 + V(23) * 3.94 + V(26) * 1 + V(27) * 1 }
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI 
M14 12 2 15 15 NMI 
G14 2 0 62 0 1m
C14  2  0 6.00P
I15 15 4 500U
V16 16 4 10.0M
GD16 16 1 TABLE { V(16,1) } ((-100,-100E-15)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -10.0M
GD13 2 13 TABLE { V(2,13) } ((-100,-100E-15)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 10.0E12
R72  2  0 10.0E12
R73  1  2 10.0E12
*C13  1  2 3.00P
*
* Noise, PSRR, and CMRR
I20 21 20 25.0
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 VALUE { 0.00 + V(3) * -28.1U + V(4) * -31.6U }
R26 26  0 1
G27  0 27 VALUE { -88.5U + V(1) * 10.0U + V(2) * 10.0U }
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 0.00
I31 0 31 DC 63.6
R31 31  0 1 TC=0.00,0.00
GD31 30 0 TABLE { V(30,31) } ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 0.00
I32 32 0 DC 85.9
R32 32  0 1 TC=0.00,0.00
GD32 0 30 TABLE { V(30,32) } ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 562M
R34  34 0 1K
C34  34 0 35.8U
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 45.4P
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 159N
E38  35 0 38 0 1
G35 33 0 TABLE { V(35,3) } ((-1,-1n)(0,0)(10.0,1n))(11.0,1))
G36 33 0 TABLE { V(35,4) } ((-11.0,-1)((-10.0,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 350
C58  5  0 2.00P
G57  0 57 VALUE { V(3) * 1.07M + V(4) * 1.42M + V(35) * 2.85M }
GD55 55 57 TABLE { V(55,57) } ((-0.2m,-1)(-0.1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE { V(57,56) } ((-0.2m,-1)(-0.1m,-1m)(0,0)(10,1n))
E55 55  0 VALUE { -325U + V(3) * 1 + V(51) * -25.0M }
E56 56  0 VALUE { 0.00 + V(4) * 1 + V(52) * -20.0M }
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE { V(50,51) } ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE { V(50,52) } ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 VALUE { -500U + V(51) * 1M }
G54  0  4 VALUE { -500U + V(52) * -1M }
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-5.10M,4.78U
G97 0 98 TABLE { V(96,5) } ((-5.6,-11.0M)(-1.00M,-10.8M)(0,0)(1.00M,10.8M)(5.6,11.0M))
E97 99 0 VALUE { V(98) * LIMIT((( V(3) - V(4) ) * 515M + -30.3M), 0.00, 1E6 ) * LIMIT((( V(3) - V(4) ) * 1.00 + -1.00), 0, 1) }
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=120U,-264N
G61 3 4 61 0 1
G60 0 61 TABLE { V(3, 4) } ((0, 0)(750M,1.08U)(1.5,100U)(2.00,100U)(3.00,102U)(5.5,108U)(6.5,120U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=2.5
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1000uA
R62 0 62 REXP  449.71912N
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1000uA
R63 0 63 REXP2  32.94705U
*
* Models
.MODEL NMI NMOS(L=2.00U W=42.0U KP=200U LEVEL=1 )
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=4.5N AF=1
.MODEL REXP  RES TCE= 5.88717
.MODEL REXP2  RES TCE= 4.7086
.ENDS MCP6471




