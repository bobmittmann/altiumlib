*
**********************************************************
*
*BCM857DS
*
* NXP Semiconductors
*
* Matched double PNP/PNP transistor
* IC   = 100 mA
* VCEO = 45 V 
* hFE  = 200 - 450 @ 5V/2mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 457
* 
* Package Pin 1;4: Emitter     	TR1;TR2
* Package Pin 2;5: Base        	TR1;TR2
* Package Pin 3;6: Collector   	TR2;TR1
*
*
* Extraction date (week/year): 47/2005
* Simulator: Spice 3
*
**********************************************************
*#
* Please note: The following model is to be used twice in 
* schematic due to equality of both transistors.
*
.SUBCKT BCM857DS 1 2 3
*
* The Diode D1, transistor Q2 and resistors RQ1 
* are dedicated to improve modeling of quasi
* saturation area and reverse mode operation
* and do not reflect physical devices.    
*
Q1 1 2 3 MAIN 0.9196 
Q2 11 2 3 MAIN 0.08035
D1 1 2 DIODE 
RQ1 1 11 111.9
*
.MODEL MAIN PNP 
+ IS = 1.619E-014 
+ NF = 0.9835 
+ ISE = 7.218E-015 
+ NE = 1.521 
+ BF = 266.9 
+ IKF = 0.08202 
+ VAF = 12.88 
+ NR = 0.977 
+ ISC = 3.672E-015 
+ NC = 1.122 
+ BR = 10.73 
+ IKR = 0.03072 
+ VAR = 24.01 
+ RB = 39.4 
+ IRB = 0.0001272 
+ RBM = 1.321 
+ RE = 0.3 
+ RC = 0.5566 
+ XTB = 0 
+ EG = 1.11 
+ XTI = 3 
+ CJE = 1.14E-011 
+ VJE = 0.7923 
+ MJE = 0.4031 
+ TF = 9E-010 
+ XTF = 20 
+ VTF = 5 
+ ITF = 0.52 
+ PTF = 0 
+ CJC = 5.839E-012 
+ VJC = 1 
+ MJC = 0.5758 
+ XCJC = 1 
+ TR = 1E-009 
+ CJS = 0 
+ VJS = 0.75 
+ MJS = 0.333 
+ FC = 0.79
*
.MODEL DIODE D 
+ IS = 5.409E-017 
+ N = 0.9852 
+ BV = 1000 
+ IBV = 0.001 
+ RS = 2.939 
+ CJO = 0 
+ VJ = 1 
+ M = 0.5 
+ FC = 0 
+ TT = 0 
+ EG = 1.11 
+ XTI = 3 
.ENDS
