*Green-Lis Macromodel Architecture
*OPAx209  Sept 3,2010 (PSpice format)
********************************************
**  This file was created by TINA      **
**    (c) 1996-2006 DesignSoft, Inc.   **
********************************************
* Rev. A by Marek Lis; Sept 3, 2010,
*
*
* This macromodel has been optimized to model the AC, DC, noise, and transient response performance within 
* the device data sheet specified limits. Correct operation of this macromodel has been verified on DesignSoft
* TINA Version 7.0.80.224 SF. For help with other analog simulation software, please consult the software supplier.
*
*  
* Copyright 2010 by Texas Instruments Corporation
* BEGIN MODEL OPA209
*GREEN-LIS MACRO-MODEL SIMULATED FEATURES:
*OPEN LOOP GAIN AND PHASE VS FREQUENCY WITH RL AND CL EFFECTS
*INPUT COMMON MODE REJECTION WITH FREQUENCY
*POWER SUPPLY REJECTION WITH FREQUENCY
*INPUT IMPEDANCE VS FREQUENCY 
*OUTPUT IMPEDANCE VS FREQUENCY
*INPUT VOLTAGE NOISE VS FREQUENCY
*INPUT CURRENT NOISE VS FREQUENCY 
*OUTPUT VOLTAGE SWING VS OUTPUT CURRENT
*SHORT-CIRCUIT OUTPUT CURRENT
*QUIESCENT CURRENT VS SUPPLY VOLTAGE
*SETTLING TIME VS CAPACITIVE LOAD
*SLEW RATE
*SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
*LARGE SIGNAL RESPONSE
*OVERLOAD RECOVERY TIME
*INPUT BIAS CURRENT
*INPUT VOLTAGE OFFSET
*INPUT COMMON MODE RANGE
*OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS
*$
.SUBCKT OPA209_0 -IN +IN V- V+ Vout
V7          40 12 -1.5
Vos         30 31 0
V11         55 56 100M
V10         57 58 100M
V6          11 63 10
V5          64 11 10
V4          60 62 12
V1          61 59 12
V9          76 13 1.5
IS2         V+ 30 0
IS1         V+ V- 2.2M
IS3         35 V- -4.5N
V3          82 11 65
V2          11 83 65
XIn11       31 32 FEMT_0
XU14        33 11 34 35 VCVS_LIMIT_0
L3          36 11 8U 
L2          37 11 1.5U 
R1          37 33 1 
GVCCS2      11 33 11 38  1
XU13        12 39 IDEAL_D_0
EVCVS5      40 11 V- 11  1
XR109       27 11 RNOISE_FREE_0
XR109_2     41 11 RNOISE_FREE_0
XR109_3     42 43 RNOISE_FREE_0
L1          43 11 75U 
C11         41 11 100P 
XR109_4     26 11 RNOISE_FREE_0
C1          11 44 63.9N IC=0 
EVCVS1      15 11 45 46  -1
R38         44 47 10 
VCCVS2_in   46 48
HCCVS2      47 11 VCCVS2_in   1K
XU9         44 11 49 50 VARICAP_0
XU7         44 11 46 51 VC_RES_0
C25         15 49 500F 
R37         50 51 26.135MEG 
C24         15 14 90N 
R32         14 49 1.8K 
R31         49 51 100MEG 
R30         15 49 500K 
EVCVS2      51 11 11 49  20MEG
GVCCS12     11 27 41 11  1M
XU5         16 11 V+ 17 VCVS_LIMIT_1
XU6         11 16 18 V- VCVS_LIMIT_1
C15         V+ V- 10P 
C22         11 23 1P
R29         23 25 1 
C23         11 28 1P 
C9          52 11 10P 
R26         52 16 10 
C21         11 19 1P 
C20         11 20 1P 
C19         21 11 1P 
C17         22 11 1P 
C16         11 53 1P 
C12         54 11 1P 
R13         45 28 1 
SW14        14 15 19 11  S_VSWITCH_1
SW13        15 14 11 20  S_VSWITCH_2
R36         28 58 1M 
R35         28 56 1M 
SW12        59 55 21 11  S_VSWITCH_3
SW11        57 60 11 22  S_VSWITCH_4
R34         28 61 1K 
R33         28 62 1K 
SW10        64 25 23 11  S_VSWITCH_5
SW9         25 63 11 23  S_VSWITCH_6
R25         65 21 1 
R19         66 22 1 
R16         67 53 1 
R14         68 54 1 
R12         69 19 1 
R7          70 20 1 
R5          71 26 10M 
R6          72 25 10M 
R4          73 24 10M 
R15         0 11 100MEG 
C13         26 11 1F 
GVCCS1      11 26 27 11  1M
GIsinking   V- 11 74 11  1M
GIsourcing  V+ 11 75 11  1M
R23         74 11 10K 
SW7         16 74 52 11  S_VSWITCH_7
R21         11 75 10K 
SW8         16 75 52 11  S_VSWITCH_8
SW4         72 69 19 11  S_VSWITCH_9
SW3         70 72 11 20  S_VSWITCH_10
XU3         60 29 70 11 VCVS_LIMIT_2
XU1         59 29 69 11 VCVS_LIMIT_2
SW2         73 65 21 11  S_VSWITCH_11
SW1         66 73 11 22  S_VSWITCH_12
XU8         30 V+ IDEAL_D_1
XU12        V- 30 IDEAL_D_1
EVCVS6      76 11 V+ 11  1
R22         77 39 100 
EVCVS4      77 11 30 11  1
XU2         39 13 IDEAL_D_0
XVn11       78 31 VNSE_0
SW6         71 67 53 11  S_VSWITCH_13
SW5         68 71 11 54  S_VSWITCH_14
XU26        39 35 11 79 VCCS_LIMIT_0
XU4         79 11 11 25 VCCS_LIMIT_1
LPSR        80 11 200M 
XVCVSPSRR   81 11 34 32 VCVS_LIMIT_3
XU22        82 16 66 11 VCVS_LIMIT_4
XU21        83 16 65 11 VCVS_LIMIT_4
XU20        18 Vout 67 11 VCVS_LIMIT_4
XU19        17 Vout 68 11 VCVS_LIMIT_5
XU11        V- 35 IDEAL_D_1
XU10        35 V+ IDEAL_D_1
C10         24 11 1F 
C5          27 11 1F
XR109_5     24 11 RNOISE_FREE_0
GVCCS15     11 24 26 11  1M
GVCCS10     11 41 42 11  1M
R20         +IN 78 100 
R18         -IN 32 100 
GVCCS6      11 42 29 11  1M
XR102       84 85 RNOISE_FREE_1
XR101       86 84 RNOISE_FREE_1
C6          84 0 1 
XR105       29 11 RNOISE_FREE_1
XR104       25 11 RNOISE_FREE_0
XR103       11 79 RNOISE_FREE_1
EVCVS34     11 0 84 0  1
C8          78 11 2P 
RPSR        80 81 1 
GVCCS11     11 81 V+ V-  50N
RCM         36 38 1 
EVCVS29     86 0 V+ 0  1
EVCVS28     85 0 V- 0  1
CinnCM      11 32 2P 
GVCCS7      11 38 30 11  350N
C7          32 78 4P 
VCCVS1_in   48 Vout
HCCVS1      16 11 VCCVS1_in   1K
GVCCS5      11 29 25 11  1U
Ccc         25 11 40U 
EVCVS3      45 11 24 11  1
.MODEL S_VSWITCH_1 VSWITCH (RON=1 ROFF=100MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1 ROFF=100MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=10MEG VON=-10M VOFF=0)
.MODEL S_VSWITCH_8 VSWITCH (RON=1M ROFF=10MEG VON=10M VOFF=0)
.MODEL S_VSWITCH_9 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_10 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_11 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_12 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_13 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_14 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.ENDS
*$
* BEGIN PROG NSE FEMTO AMP/RT-HZ 
.SUBCKT FEMT_0  1 2
* BEGIN SETUP OF NOISE GEN - FEMPTOAMPS/RT-HZ
* INPUT THREE VARIABLES
* SET UP INSE 1/F
* FA/RHZ AT 1/F FREQ
.PARAM NLFF=3.8E3
* FREQ FOR 1/F VAL
.PARAM FLWF=.1
* SET UP INSE FB
* FA/RHZ FLATBAND
.PARAM NVRF=500
* END USER INPUT
* START CALC VALS
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
*$
* END PROG NSE FEMTO AMP/RT-HZ
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS 
*$
*TG IDEAL DIODE
.SUBCKT IDEAL_D_0  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS
*$
* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS 
*$
*VARICAP (VOLTAGE-CONTROLLED CAPACITOR
.SUBCKT VARICAP_0  1 2 3 4
*PINS       VC+ VC- CAP+ CAP-
R1 3 10 1U
VC 10 20 0
EC 20 4 VALUE = {(1/(((ABS(V(1,2))*(-2.08)+104.636))))*V(INT)*100000000000000000}
GINT 0 INT VALUE = {I(VC)}
CINT INT 0 1
RINT INT 0 10e6
.ENDS
*$
*VOLTAGE CONTROLLED RESISTOR
.SUBCKT VC_RES_0  1      2      3    4
*              VC+    VC-   RES1 RES2
ERES 3 40 VALUE = {(I(VSENSE) * (ABS(V(1,2))*ABS(V(1,2))*0.000352-0.02359*ABS(V(1,2))+0.5922))*140000*24200*50*2/414500}
VSENSE 40 4 DC 0
.ENDS
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VC+ VC- VOUT+ VOUT-
*              
E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = (0,0.2) (30,0.6) (50,1.5) (64, 2.5)
.ENDS 
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 6000
.PARAM VNEG = -6000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS
*$
*TG IDEAL DIODE
.SUBCKT IDEAL_D_1  A C
D1 A C DNOM 
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS
*$
* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=1
* FREQ FOR 1/F VAL
.PARAM FLW=50
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=0.25
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
*$
* END PROG NSE NANOV/RT-HZ
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 1M
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),IPOS,INEG)}
.ENDS
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_1  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 6
.PARAM IPOS = 250
.PARAM INEG = -250
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),IPOS,INEG)}
.ENDS
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_3  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = -1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_4  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS
*$
*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_5  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VPOS,VNEG)}
.ENDS
*$
* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS
.END
*$
