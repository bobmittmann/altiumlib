*Rev.a May-2007
* BEGIN MODEL LMV551
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THRU
* THE SUPPLY RAILS, OUTPUT SWING VS IO, OUTPUT CURRENT LIMIT,
* OPEN LOOP GAIN AND PHASE, SLEW RATE, COMMON MODE REJECTION
* WITH FREQ EFFECTS, POWER SUPPLY REJECTION WITH FREQ EFFECTS,
* INPUT VOLTAGE NOISE WITH 1/F, INPUT CURRENT NOISE WITH 1/F,
* INPUT CAPACITANCE, INPUT BIAS CURRENT VS TEMPERATURE, INPUT
* COMMON MODE RANGE, INPUT OFFSET VS TEMPERATURE, HIGH CLOAD
* EFFECTS, AND QUIESCENT CURRENT VS VOLTAGE AND TEMPERATURE.
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  1   3   5  2  4
.SUBCKT LMV551 1 3 5 2 4
Q20 6 7 8 QLN
R3 9 10 2E3
R4 9 11 2E3
R10 7 12 1E3
R11 13 14 1E3
R12 15 5 8
R13 2 16 8
R16 17 18 10E3
R17 19 20 8
R18 8 21 8
D5 4 5 DD
D6 2 4 DD
D7 22 0 DIN
D8 23 0 DIN
I8 0 22 0.1E-3
I9 0 23 0.1E-3
E2 8 0 2 0 1
E3 20 0 5 0 1
D9 24 0 DVN
D10 25 0 DVN
I10 0 24 1E-3
I11 0 25 1E-3
E4 26 3 24 25 19E-3
G2 27 3 22 23 3E-6
R22 2 5 5E6
E5 28 0 20 0 1
E6 29 0 8 0 1
E7 30 0 31 0 1
R30 28 32 1E5
R31 29 33 1E5
R32 30 34 1E5
R33 0 32 10
R34 0 33 10
R35 0 34 10
E10 35 1 34 0 3E-2
R36 36 31 1E3
R37 31 37 1E3
C6 28 32 1E-12
C7 29 33 1E-12
C8 30 34 1E-12
E11 38 35 33 0 0.2
E12 27 38 32 0 -0.48
E14 39 8 20 8 0.6
D11 17 20 DD
D12 8 17 DD
M1 40 41 16 16 NOUT L=3U W=400U
M2 42 43 15 15 POUT L=3U W=400U
M3 44 44 19 19 POUT L=3U W=400U
M8 45 45 21 21 NOUT L=3U W=400U
R43 46 43 100
R44 47 41 100
G3 17 39 48 39 0.125E-3
R45 39 17 9.2E6
C12 18 49 3.6E-12
R46 50 51 2
R47 52 51 2
C13 10 11 2E-12
C14 27 0 1E-12
C15 26 0 1E-12
C16 4 0 3E-12
D13 41 6 DD
D14 53 43 DD
Q15 53 14 20 QLP
V18 54 55 0.8E-3
E17 37 0 27 0 1
E18 36 0 3 0 1
V21 9 8 0
R59 56 42 40
R60 40 57 10
J1 58 27 58 JNC
J2 58 26 58 JNC
J3 26 59 26 JNC
J4 27 59 27 JNC
E20 60 39 11 10 1
R62 60 48 1E4
C23 48 39 4E-12
G7 61 39 17 39 -1E-3
G8 39 62 17 39 1E-3
G9 39 63 45 8 1E-3
G10 64 39 20 44 1E-3
D17 64 61 DD
D18 62 63 DD
R66 61 64 100E6
R67 63 62 100E6
R68 64 20 1E3
R69 8 63 1E3
E23 20 46 20 64 1
E24 47 8 63 8 1
R70 62 39 1E6
R71 63 39 1E6
R72 39 64 1E6
R73 39 61 1E6
R75 38 27 1E9
R76 35 38 1E9
R77 1 35 1E9
R78 3 26 1E9
R79 39 48 1E9
R81 46 20 1E9
R82 8 47 1E9
R83 31 0 1E9
G14 65 8 66 0 15.37E-6
G15 44 45 66 0 15E-6
V51 66 0 1
I21 5 2 18.5E-6
V78 20 58 0
V79 59 8 0.2
R155 44 20 1E8
R156 8 45 1E8
R157 16 41 1E8
R158 15 43 1E8
E98 20 13 5 15 8
E99 12 8 16 2 3.5
R336 17 49 5.5E8
R340 0 66 1E12
R341 0 66 1E12
R342 55 67 127K
R343 26 68 127K
E100 49 0 4 0 1
I22 27 0 19E-9
I23 26 0 19E-9
G25 27 3 69 70 3.7E-6
R409 0 69 5E4
R410 0 69 5E4
R411 0 70 5E4
R412 0 70 5E4
V127 56 4 0.070
V128 4 57 0.125
I31 0 71 1E-3
D31 71 0 DD
R415 0 71 1E9
V131 71 72 0.65
R416 0 72 2E9
G26 5 2 72 0 -6E-5
G27 27 0 72 0 -2E-8
G28 26 0 72 0 -2E-8
E120 27 54 72 0 3.3E-3
V133 73 51 0.09
M21 10 67 52 52 PIN L=3U W=90U
M22 11 68 50 50 PIN L=3U W=90U
M23 65 65 20 20 PIN L=3U W=90U
M24 73 65 20 20 PIN L=3U W=90U
R418 65 20 1E12
R419 0 72 2E9
C35 54 0 1E-15
.MODEL DVN D KF=9E-12 IS=1E-16
.MODEL DD D
.MODEL DIN D KF=9E-16 IS=1E-16
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL JNC NJF IS=1E-18
.MODEL POUT PMOS KP=200U VTO=-0.7
.MODEL NOUT NMOS KP=200U VTO=0.7
.MODEL PIN PMOS KP=200U VTO=-0.7
.ENDS
* END MODEL LMV551
