* MAX4714 MACROMODEL
* ------------------------------
* Revision 0, 10/2004
* ------------------------------
* MAX4714 is a low-voltage, low on-resistance, single single-pole/double throw
* analog switch operating from a single +1.6V to +3.6V supply.
* ------------------------------
* Connections
*      1  = IN
*      2  = V+
*      3  = GND
*      4  = NC 
*      5  = COM
*      6  = NO
*****************
.SUBCKT MAX4714 1 2 3 4 5 6
X1 6 4 5 1 2 3 MAX4714SPDT
.ENDS
*****************
***************** 
.SUBCKT MAX4714SPDT 1 2 3 4 5 6 
S1 1 3 4 6 SMOD1
S2 2 3 4 6 SMOD2
*SUPPLY CURRENT
RSUPP 5 3 90MEG
*ANALOG SIGNAL RANGES
DCOM1 3 5 DX
DCOM2 6 3 DX
DNO1 1 5 DX
DNO2 6 1 DX
DNC1 2 5 DX
DNC2 6 2 DX
*CHARGE-INJECTION
CNOIN 4 1 23.5P
CNCIN 4 2 23.5P
CCOMIN 4 3 23.5P 
*FREQUENCY RESPONSE OF OFF-ISOLATION
CNOI 1 3 5.65P
CNCI 2 3 5.65P
*ON/OFF-CAPACITANCE
ELOGIC 16 6 4 6 1
DLH 16 17 DX
DLL 18 16 DX
VLH 17 19 1.4 
VLL 18 19 0.5
RSC 19 20 1
VIMEAS 20 6 0
FDIS 6 21 VIMEAS 1
DL 6 21 DX
DH 21 22 DX
VCLAMP 22 6 1
RPU 21 23 1MEG
VPU 23 6 0.5
GSCALED 6 24 21 6 1
VSCALED 24 6 0
FDISI 27 6 VIMEAS 1
DLI 6 27 DX
DHI 27 28 DX
VCLAMPI 28 6 1
RPUI 27 29 1MEG
VPUI 29 6 0.5
GSCALEDI 6 30 27 6 1
VSCALEDI 30 6 0
**
CNOT 1 25 1.45P
VNOT 25 6 0
FNOT 1 6 POLY(2) VNOT VSCALED 0 0 0 0 8.05
**
CNCT 2 26 1.45P
VNCT 26 6 0
FNCT 2 6 POLY(2) VNCT VSCALEDI 0 0 0 0 8.05
*MODELS USED
.MODEL SMOD1 VSWITCH(RON=0.6 ROFF=62.946E6 VON=1.4 VOFF=0.5)
.MODEL SMOD2 VSWITCH(RON=0.6 ROFF=62.946E6 VON=0.5 VOFF=1.4)
.MODEL DX D(IS=1E-18 N=0.001)
.ENDS
*****************

* Copyright (c) 2003-2012 Maxim Integrated Products.  All Rights Reserved.
