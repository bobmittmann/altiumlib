**************** Power Discrete MOSFET Electrical Circuit Model *****************
* Product Name: FQT5P10
* 100V P-Channel MOSFET and SOT-223
*--------------------------------------------------------------------------------
.SUBCKT FQT5P10 20 10 30
Rg 10 1  0.077
M1 2 1 3 3 DMOS  L=1u  W=1u
.MODEL DMOS PMOS (VTO={-3.8*{-0.0005*TEMP+1.0125}} KP={2.45*{-0.00002*TEMP+1.0005}}
+ THETA=0.0576  VMAX=1.0E5   LEVEL=3)
Cgs 1 3 240p
Rd 20 4 0.273  TC=0.0081
Dds 4 3 DDS
.MODEL DDS D(BV={100*{0.000875*TEMP+0.978125}}  M=0.37   CJO=52p   VJ=0.609)
Dbody 20 3 DBODY
.MODEL DBODY D(IS=1.0E-14  N=1.0  RS=0.34  EG=1.18  TT=85n)
Ra 4 2  0.273  TC=0.0081
Rs 3 5  0.022
Ls 5 30 2.6n
M2 1 8 6 6 INTER
E2 8 6 4 1 2
.MODEL INTER PMOS (VTO=0 KP=10 LEVEL=1)
Cgdmax 7 4 380p
Rcgd 7 4 1E7
Dgd  4 6 DGD
Rdgd 4 6 1E7
.MODEL DGD D(M=0.77 CJO=380p VJ=0.44)
M3 7 9 1 1 INTER
E3 9 1 4 1 -2
.ENDS
*-------------------------------------------------------------------------------
* Creation : Feb.-14-2005
* Fairchild Semiconducto

