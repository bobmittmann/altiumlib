* BEGIN MODEL LM7321
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*///////////////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   4   5  2  1
.SUBCKT LM7321 3 4 5 2 1
* SEE BELOW FOR PROGRAMMING INFORMATION
* SEE BELOW FOR MODEL FEATURES
* START PROGRAMMING
* BECAUSE THE PARAMETERS OF THE LM7321 VARY NOTICABLY AND NONLINEARLY
* WITH OPERATING VOLTAGE OVER THE WIDE OPERATING VOLTAGE RANGE OF THE
* PART (2.7 TO 30 VOLTS), THE MODEL IS PROGRAMMABLE TO SOME EXTENT.
* THERE ARE THREE GROUPS OF SPICE STATEMENTS FOR PROGRAMMING. ONLY
* ONE GROUP SHOULD BE UN-COMMENTED AT A TIME. THE THREE GROUPS ARE
* FOR 2.7, 10, AND 30 VOLTS TOTAL ACROSS THE PART. THE MODEL IS NOW
* SET UP FOR 30 VOLTS IE THE 30 VOLT GROUP IS UN-COMMENTED. FOR OTHER
* SUPPLY VOLTAGES THE VALUES MAY BE INTERPOLATED. SEE BELOW FOR AN
* INDEX TO THE FUNCTIONS OF THE PROGRAMMABLE COMPONENTS. V6 AND V7
* MAY BE ADJUSTED FOR ANY DESIRED OFFSET OR OFFSET DELTA FOR INPUT
* COMMON MODE NEAR THE POSITIVE RAIL. NOTE THAT BECAUSE THE MODEL
* HAS REALISTIC COMMON MODE AND POWER SUPPLY REJECTION, THE OFFSET
* WILL CHANGE WITH SUPPLY VOLTAGES AND COMMON MODE VOLTAGE.
*
* 30 VOLT TOTAL SUPPLY GROUP
C24 16 28 5.6E-12
R159 20 15 2E6
R219 15 28 8E7
R316 47 44 60
R317 47 46 60
R318 54 59 60
R319 51 59 60
R320 60 61 4.4E3
R324 65 45 4.4E3
I16 5 2 1.33E-3
G25 5 2 42 0 -3.3E-3
F1 5 2 V15 -0.23
R153 15 16 500
E152 82 81 75 0 0.37
C29 71 75 150E-12
E151 81 78 76 0 -0.53
V6 43 53 -600E-6
V7 61 53 2.7E-3
E158 60 82 42 0 1.125E-3
E150 78 3 77 0 3.3E-3
E84 13 10 13 12 6.0
E85 9 8 14 8 3.65
E146 65 70 68 69 0.6
G30 60 65 89 0 8E-5
G27 60 65 66 67 1.7E-4
* END 30 V TOTAL SUPPLY GROUP
*
* 10 VOLT TOTAL SUPPLY GROUP
*C24 16 28 8.2E-12
*R159 20 15 1.2E6
*R219 15 28 3E7
*R316 47 44 55
*R317 47 46 55
*R318 54 59 55
*R319 51 59 55
*R320 60 61 5.3E3
*R324 65 45 5.3E3
*I16 5 2 1.1E-3
*G25 5 2 42 0 -2.5E-3
*F1 5 2 V15 -0.12
*R153 15 16 400
*E152 82 81 75 0 0.22
*C29 71 75 150E-12
*E151 81 78 76 0 -0.75
*V6 43 53 -600E-6
*V7 61 53 2.0E-3
*E158 60 82 42 0 1.125E-3
*E150 78 3 77 0 2E-3
*E84 13 10 13 12 4.6
*E85 9 8 14 8 3.75
*E146 65 70 68 69 0.6
*G30 60 65 89 0 8E-5
*G27 60 65 66 67 1.7E-4
* END 10 V TOTAL SUPPLY GROUP
*
* 2.7 VOLT TOTAL SUPPLY GROUP
*C24 16 28 11.5E-12
*R159 20 15 5E5
*R219 15 28 1.3E7
*R316 47 44 42
*R317 47 46 42
*R318 54 59 42
*R319 51 59 42
*R320 60 61 3.6E3
*R324 65 45 3.6E3
*I16 5 2 1.1E-3
*G25 5 2 42 0 -3.3E-3
*F1 5 2 V15 -0.12
*R153 15 16 500
*E152 82 81 75 0 -0.57
*C29 71 75 1E-12
*E151 81 78 76 0 0.42
*V6 43 53 -350E-6
*V7 61 53 1.2E-3
*E158 60 82 42 0 8.8E-4
*E150 78 3 77 0 -1E-3
*E84 13 10 13 12 6.3
*E85 9 8 14 8 4.6
*E146 65 70 68 69 0.55
*G30 60 65 89 0 8E-6
*G27 60 65 66 67 6.9E-5
* END 2.7 V TOTAL SUPPLY GROUP
*
* END PROGRAMMING
* INDEX TO SOME PROGRAMMABLE COMPONENT FUNCTIONS
* THE LINES IN THIS INDEX MUST ALWAYS REMAIN COMMENTED
*
*V6    RELATIVE OFFSET BETWEEN INPUT STAGES
*V7    OVERALL  OFFSET
*E158  TEMCO OF OFFSET
*
* END OF INDEX
*
* MODEL FEATURES INCLUDE GAIN AND PHASE, SLEW RATE,
* VOLTAGE NOISE WITH 1/F, CURRENT NOISE WITH 1/F,
* INPUT BIAS CURRENT, INPUT BIAS CURRENT CHANGE
* WHEN COMMON MODE VOLTAGE NEAR THE + RAIL, INPUT
* OFFSET VOLTAGE, INPUT OFFSET VOLTAGE CHANGE WHEN
* WHEN COMMON MODE VOLTAGE NEAR THE + RAIL, INPUT
* OFFSET TEMPCO, COMMON MODE RANGE, CMRR WITH FREQ
* EFFECTS, PSRR WITH FREQ EFFECTS, OUTPUT SWING,
* OUTPUT CURRENT FLOWS THROUGH THE RAILS, OUTPUT
* CURRENT LIMIT, IQ, IQ TEMPCO, AND IQ CHANGE WITH
* COMMON MODE VOLTAGE, AND CAPACATIVE LOAD EFFECTS.
*
Q41 6 7 8 QLN
R148 7 9 1E3
R149 10 11 1E3
R150 12 13 2.7
R151 8 14 2.7
R154 17 13 2.7
R155 8 18 2.7
D22 19 5 DD
D23 2 19 DD
E58 8 0 2 0 1
E79 13 0 5 0 1
R156 2 5 1.1E5
E60 20 8 13 8 0.5
D24 21 13 DD
D25 8 22 DD
R157 23 24 100
R158 25 26 100
G14 15 20 27 20 0.1E-3
C25 19 0 0.5E-12
D26 26 6 DD
D27 29 24 DD
Q42 29 11 13 QLP
R160 19 30 1
R161 31 19 1
E71 32 20 33 34 -1
R162 32 27 1E3
C26 27 20 0.1E-12
G15 35 20 15 20 -1E-3
G16 20 36 15 20 1E-3
G17 20 37 38 8 1E-3
G18 39 20 13 40 1E-3
D28 39 35 DD
D29 36 37 DD
R163 35 39 1E9
R164 37 36 1E9
R165 39 13 1E3
R166 8 37 1E3
R167 36 20 1E7
R168 37 20 1E7
R169 20 39 1E7
R170 20 35 1E7
R171 20 27 1E9
R172 23 13 1E9
R173 8 25 1E9
G20 40 38 41 0 90E-6
L2 19 1 0.4E-9
R175 19 1 4E2
R176 40 13 1E8
R177 8 38 1E8
R178 14 26 1E8
R179 12 24 1E8
E24 28 0 19 0 1
Q52 30 24 12 QOP
Q53 31 26 14 QON
Q54 38 38 18 QON
Q55 40 40 17 QOP
E144 13 23 13 39 1
E145 25 8 37 8 1
E51 15 22 20 8 0.9
E52 21 15 13 20 0.9
G23 5 0 30 19 1
G24 2 0 19 31 -1
Q56 33 43 44 QIN
Q57 34 45 46 QIN
Q58 47 48 8 QLN
Q59 48 49 8 QLN
Q60 50 45 51 QIP
Q61 52 53 54 QIP
Q62 55 56 13 QLP
Q63 48 57 58 QPX
R321 33 62 350
R322 63 50 350
R323 63 52 350
V4 13 64 1
D30 43 13 DD
D31 45 13 DD
D32 8 53 DD
D33 8 45 DD
D34 66 0 DIN
D35 67 0 DIN
I9 0 66 0.1E-3
I10 0 67 0.1E-3
C27 60 0 1E-12
C28 4 0 1E-12
D36 68 0 DVN
D37 69 0 DVN
I11 0 68 0.1E-3
I12 0 69 0.1E-3
E147 71 0 13 0 1
E148 72 0 8 0 1
E149 73 0 74 0 1
R329 71 75 1E6
R330 72 76 1E6
R331 73 77 1E6
R332 0 75 100
R333 0 76 100
R334 0 77 1E4
R335 79 74 1E3
R336 74 80 1E3
C30 72 76 1E-12
C31 73 77 1E-12
R337 34 62 350
C32 34 33 2E-12
C33 50 52 2E-12
G28 15 20 83 20 0.1E-3
E153 84 20 50 52 1
R338 84 83 1E3
C34 83 20 0.1E-12
R339 20 83 1E9
V12 41 0 1
V15 55 59 0
R341 55 58 1
R342 57 64 1
R343 48 49 8E-2
I14 0 85 1E-3
D39 85 0 DD
R345 0 86 1E7
E155 87 0 86 0 -1.75
R346 0 87 1E7
V17 85 86 1.2301
G29 13 56 87 0 -30E-6
E156 70 4 88 0 1.25E-6
R347 0 88 9.6E4
R348 0 88 9.6E4
R349 0 89 1E4
R350 0 89 1E4
I15 0 90 1E-3
D40 90 0 DD
R352 0 42 1E7
V19 90 42 0.655
R353 82 60 1E9
R354 81 82 1E9
R355 78 81 1E9
R356 3 78 1E9
R357 0 41 1E9
E159 80 0 60 0 1
E160 79 0 65 0 1
V21 13 62 -0.3
V22 63 8 -0.3
.MODEL QON NPN RC=1 IS=1E-13
.MODEL QOP PNP RC=1 IS=1E-13
.MODEL QPX PNP BF=200 IS=1E-14
.MODEL DD D
.MODEL QIN NPN BF=3200
.MODEL QIP PNP BF=1350
.MODEL DVN D KF=2.5E-15
.MODEL DIN D KF=1E-15
.MODEL QLN NPN
.MODEL QLP PNP
.ENDS
* END MODEL LM7321
