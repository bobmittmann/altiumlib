*SRC=DMP2066LDM;DI_DMP2066LDM;MOSFETs P;Enh;20.0V 4.60A 40.0mohms
*SYM=POWMOSP
.SUBCKT DI_DMP2066LDM   10 20 30
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  18.0m
RS  40  3  2.00m
RG  20  2  32.6
CGS  2  3  660p
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.47n
R1  13  0  1.00
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1.00
D2  15  0  DLIM
DSD  10 3  DSUB
LS  30 40  7.50n
.MODEL DMOS PMOS(LEVEL=3 VMAX=41.7k THETA=80.0m
+ ETA=2.00m VTO=-1.20 KP=43.8
.MODEL DCGD D (CJO=1.47n VJ=0.600 M=0.680
.MODEL DSUB D (IS=19.1n N=1.50 RS=0.141 BV=20.0
+ CJO=350p VJ=0.800 M=0.420 TT=223n
.MODEL DLIM D (IS=100U)
.ENDS
