**$ENCRYPTED_LIB
**$INTERFACE
*****************************************************************************
* (C) Copyright 2013 Texas Instruments Incorporated. All rights reserved.
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer.
*****************************************************************************
*
** Released by: WEBENCH(R) Design Center, Texas Instruments Inc.
* Part: SN74VC2G66_Q1
* Date: 06/25/2013
* Model Type: All In One
* Simulator: PSPICE
* Simulator Version: 16.2.0.p001
* EVM Order Number: N/A
* EVM Users Guide: N/A
* Datasheet: SCES829A
* 
* Model Version: 1.0
* 
*****************************************************************************
* 
* Updates: 
* 
* Version 1.0 : Release to Web
* 
*****************************************************************************
* 
* Notes:The following will be modeled for 4.5V supply :
*VIH, VIL, VI/O, Ron, IS(off), IS(on), Ii(control input current), 
*ICC, Cic, Cio(off) Cio(on), ten=tdis, frequency response and sinewave distortion
*****************************************************************************

.SUBCKT SN74VC2GG66_Q1 A GND C B VDD
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
bd5b78ae38739119cb47925e363f50c5efd156fbcd784a4f197b36855ab218f42a8a2bfd4fe2703eaf193f1b96e24aebd84deecc57bef0f5a0af6402bc9c566d
12d2018c778dc7a58d95be0fc5d68720c31e684d4b0dafc804fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e5442b05feec11b7426dc8bf56258e28b
36ec8c7d9856573290c9c14c58835e14db6e6e6353859eceb1f9f3d89ff16ce77045c65ddb608a2c76b807b1a1c84e6a9e4e6f45fdc37acb12dfcc2655d11e0e
6f4f6f21b39202b4c876379922ed059f0b2654cc8404a7e829ea36acf14f2335dc78019e6b0a9af3eed94a205c1e424df1306b3e07b3eddbe3adbed052508a42
45f4bb15bdf6921e7661689f22f7c81e0bf566ccb86d9f7e93948ed3da14781e46c907e75ffa80f2197b36855ab218f42a8a2bfd4fe2703e8767c7dd05e0f608
0ab3eab7d19021d29b950a87f5202e0a6b84e67425011d333e0ccf12ae42c6862d217c8c0391442804fc163d1408fe336c2f314c02bd115cfdf5ee4f02f369e5
e8a3dc121b162709b7b7a9e62a826ce4155ee0085d73d04a93948ed3da14781e46c907e75ffa80f2197b36855ab218f42a8a2bfd4fe2703e8767c7dd05e0f608
e175e46269ccd732889d292989282f322b64ed5f6218fa888a9f10b7655494f58ade6ebda763938c01c1bb9f962af3b1afd42b708595ddfd22d51deb16fdb32d
6bfb5d61ac69ca8fc440270b84182547a26f66e77ed41af48a9f10b7655494f58ade6ebda763938c01c1bb9f962af3b1afd42b708595ddfd22d51deb16fdb32d
c36f86d7f8415e318d95be0fc5d68720989fa906b6b88ed1eed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823
8548215614db6af375d633cacd9ba862303d7240d8c3139d197b36855ab218f42a8a2bfd4fe2703eaf193f1b96e24aebd84deecc57bef0f5a0af6402bc9c566d
a0e938c77ef85915cb47925e363f50c5c6e28a73ab7cb8b604fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e5442b05feec11b7426dc8bf56258e28b
bf6e10e5e4a954b2671480172c6f865875def76a9d391d2b48d802109cddcc50eed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628ac37857e2170d31c
d1eef0ba38bb40388d95be0fc5d68720219ec249b6ed8bbad91a973676d20455e847dda77d5f9443c92c652c5889c7dfaedffb309d4ac06d35de757aa34a29ed
f6ac43e363a110959f9754c4f2799f95790b803f4746c90ec3957dac49f48ddd96898b04fbbfb16d74987d5ef2f6c63a95918ac700906ea3155f4c22fc09ee2c
274f7c635cc50221ef725d869070d679374fb235878b195aa863bd2c702c625109c3ffe26adc1589c3957dac49f48ddd96898b04fbbfb16dd84225fb11e810be
83d256eb2b3ed6e6b17f03b65f46c771bc0f55aa2a7c7b9ff3afd7464215d3049bdf9e0525a59fd2afd42b708595ddfdab66c0c1f04149e2cbc379236612eefc
8b4937c63a589ad389521aea768f7f20374fb235878b195aa863bd2c702c6251d07114f87278901ec3957dac49f48ddd96898b04fbbfb16dd84225fb11e810be
227fab7dacf394793ddd4f4aa6d81617bc0f55aa2a7c7b9ff3afd7464215d3042928868d9d3eea79afd42b708595ddfdab66c0c1f04149e2cbc379236612eefc
c466d030111bc2faf5fe1e846882b4ac6e663b4de9531360127b390fff4107f7f339d803c60d5c4ccf175441f5661e6fdbe86c1f70c2d0d34e43d4650fa78566
42ab3a9c368d14ffb9d1f2f687d0a533f96bce6ec923602e2f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
42ab3a9c368d14ffb9d1f2f687d0a5333cf74c17f52858ce2f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
42ab3a9c368d14ffb9d1f2f687d0a533bb346e603773c3ae2f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
42ab3a9c368d14ffb9d1f2f687d0a533e6b838048f27b3a92f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
$CDNENCFINISH
.ENDS

.SUBCKT SN74VC2G66_Sch_0 A GND B CNTL
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
bd5b78ae38739119f73e1ed7b8ea4c1dcc3a724096abf9f204fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e5442b05feec11b7426dc8bf56258e28b
6bfb5d61ac69ca8fe43c2769e3124dadff738c9aeff0e882c315775dd3cb52f604fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e835710869e931e5d
a978e94c36773adb8a07603bbd943ff4cdee2c5d1ef02a3e245bb2f8cad0f0d639800334b527cca10575648ea034995dafd42b708595ddfd22d51deb16fdb32d
282c5c516cd64a8c761c50ae52f536db328bc67db2e43b8b9fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5fc95b8965c803077a
2fe921c25199d9b2761c50ae52f536db7a36bfc1c891b6c6eed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823
e60c944eb0265a2521503cc3350af00b5cb58db196c68e6ceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823
7ab0454a9d7ac522ba78e90b8b71bcb18522e2b2f6352a7ba863bd2c702c625109c3ffe26adc1589c3957dac49f48ddd96898b04fbbfb16dd84225fb11e810be
07d517d38b0949d4593822f2d9e81979204f1448b85104619fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5fc95b8965c803077a
a7d0050396c3b12d6467a481ccc56229c77598dc460100a53e199232fb035d5d6a0efa8cffb1c72beed94a205c1e424df1306b3e07b3eddbe3adbed052508a42
83d256eb2b3ed6e677a6b5714f195acd8522e2b2f6352a7ba863bd2c702c6251d07114f87278901ec3957dac49f48ddd96898b04fbbfb16dd84225fb11e810be
48e1e9459b017b0ae0f086af9e9a7668e1cb4fa691e6e0e38ded7c79edb562c39fb942d9716e294013179c8d01115b803988149c093b18571396f67a589400b2
65938c97d4f143a510caf7e5a8a29a1da55e741cba0e97213a101d8231a0c597c3957dac49f48ddd96898b04fbbfb16d74987d5ef2f6c63a5ecb9e4307d35de3
36ec8c7d9856573290c9c14c58835e14db6e6e6353859eceb1f9f3d89ff16ce7c29f0c99abb8b6c42f42acd636f67afeb5bfbe0382509d5b0c09033e92d625f7
73e1090e429f354ce9ad93d47d651a3c6ed82fc3d7cf1cfd9fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5fc95b8965c803077a
c36f86d7f8415e31e9ad93d47d651a3c121b2e3708880dcceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823
e433ed7472ee6dd3e0f086af9e9a7668be5ead5c0ec814cdcdf83ffd856ffcceeed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628ac37857e2170d31c
8cc5b1271dd8a4246d227265d6691f4a9c0ba7ceb1c4dd1e1801f442a050c66e04fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e835710869e931e5d
85551fcb960525bf17d9aa03d68d78fcc77598dc460100a53e199232fb035d5dbbfc6111f3fa81efeed94a205c1e424df1306b3e07b3eddbe3adbed052508a42
35b9107f8ed5e5a5de997b41e018a6c574ed732edaed1adceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823
274f7c635cc502219f9a889e2c1ab2728522e2b2f6352a7ba863bd2c702c6251d0c5f6593ec4e0a3c3957dac49f48ddd96898b04fbbfb16dd84225fb11e810be
5ea0817094e0792a47aa5db31001657d48050618c5d4dc0d9fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5fc95b8965c803077a
c466d030111bc2faf5fe1e846882b4ac6e663b4de9531360127b390fff4107f75749fba4ad342944402fcf20637538fbdbe86c1f70c2d0d34e43d4650fa78566
d7072740a938f0e77ebf0621ad1c8d79f170c2cee7c6dbfe87292f321b3ce12f4b2136dbcfb0192c434cda99534fc92de53b26cf6c1207b580b0d1da1390d472
bf921d7c43347b936d7c83cdd3f4c7454615839ab8739af9de54eaaef8c1f9c513cc30dac1759566647a420e9970e9f1644126c9831a96bd1ebb60e3d1b7c7ba
0f65e6141a24ff98bf017e60635b36dce3362d053423d73d117e5c19a0de9911dbe86c1f70c2d0d3d22f36355734485498459f8d9427cf6d749fb528e856a8df
42ab3a9c368d14ffb9d1f2f687d0a533f96bce6ec923602e2f0ffddeaf2b0c71e80c861f82692b92c1846234f9d070371a917ca1e1150551bf970eb4406f3147
42ab3a9c368d14ffb9d1f2f687d0a5333cf74c17f52858ce2f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
42ab3a9c368d14ffb9d1f2f687d0a533bb346e603773c3ae2f0ffddeaf2b0c71f314e6fbc5b80613cf87980ba39c3f1c2bb4ba6267ec34a776c03a7ef54c51e0
42ab3a9c368d14ffb9d1f2f687d0a533e6b838048f27b3a92f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
42ab3a9c368d14ffb9d1f2f687d0a53368e3d3b6ef1a42f52f0ffddeaf2b0c71e80c861f82692b92f50e5b1b63302cd333386b78bea576bbd38aff4e12555a5d
$CDNENCFINISH
.ENDS



**** 2 INPUT AND **********************************
.SUBCKT AN210_0  A B Y DVDD DVSS PARAMS: RDRV=10K RDLY=10K CDLY=0.1PF DIV=2
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
79e116ed52a7f63d317f2b4afb6de79ceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55d65d71c5856906f8a793e969bbc00e471
e1d4d034569ddb59f3cba33b6c977327dbe86c1f70c2d0d3d22f36355734485498459f8d9427cf6dbfb94d64dccce65cb425cc4f9b2e15f453d44eb387efa1e0
d66c2b6cf650a2e3317f2b4afb6de79ceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55d65d71c5856906f8a793e969bbc00e471
764eab282c403481f3cba33b6c977327dbe86c1f70c2d0d3d22f36355734485498459f8d9427cf6dbfb94d64dccce65cb425cc4f9b2e15f453d44eb387efa1e0
f5b0f0bb8c25915b28f84a1a2d7ca963ee1fcbe4e88889f8b45fb555070e0f5886c7072f904ece1785758e5130d42cf396cd4d6b9e1c4fc489c2f78cd5fd82be
9ed557ec13469cd31cde7e44b5902cf6a0b9ff23883894aba2827a20f24dfec0dbabfd65cbdea9d4be2108b728a7f10404fc163d1408fe3330be4810d52f68d8
55d7fa3e9be65c06164eddddf70b2d309fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5f6ae4ebc7ec1b256e8f1dcd694cbf6acb
b0fb583fca8a2e0160807eda7bc0b4c3e71f71e187584171c92c652c5889c7dfaedffb309d4ac06d2c744c4029838b320afdd7f44b471c71fca3a0227cb74238
1dedaa6f0a7bf456d9ab01cc66173203bfcc361f37c6b28b9fb942d9716e294013179c8d01115b803988149c093b185760e124bd65f6dd5fc95b8965c803077a
0111d96991417d236131abc31f305113dbe86c1f70c2d0d3d22f36355734485498459f8d9427cf6dbfb94d64dccce65cb425cc4f9b2e15f453d44eb387efa1e0
5a10a0e5d71a9276317f2b4afb6de79ceed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55d65d71c5856906f8a793e969bbc00e471
$CDNENCFINISH
.ENDS AN210_0  


.SUBCKT 2TO1MUX_0  V1 V2  A  OUT    PARAMS:  VTHRESH=0.5 
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
adc2f33f705d234bea3cc43f69f7f53cdc051b9a91e3562feddd8e3ca8357da21b4fb3137ccec2da2e0dfac773813e22231d328f694806619b4a12e5afaac291
$CDNENCFINISH
.ENDS 2TO1MUX_0 




.SUBCKT VI_HL_0  VIN VDD VOUT 

$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
c0a34efabb889ecb8d5b93a323f7ddf9ecd79bd44dcc3ec33a948fb397a15d052bce9f27643691805f3b65bef6c937658184edbb04a995fed38aff4e12555a5d
55c1fc83d899a54353ff0e45f24888d3782abd8ef87334bb93679504deb73bcd9c6d52ccecb6cab4b77d9a0e757baf9cafd42b708595ddfd22d51deb16fdb32d


$CDNENCFINISH
.ENDS  



.SUBCKT COMP_0  VDD VP VN VO VSS

*///////////////////////////////
*//
*// BEGINS MODEL
*//

$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
e93c5c830b64d2dbd9b337e692a73b4372957c6cd8e026764a04a731b09ab3f8c481d5b1c27c2d50be2108b728a7f10404fc163d1408fe3330be4810d52f68d8
0ef271de5a0e4e2a41c641296792e5d32d1975fe69f1273ee2af75b8445acede59ceb4be71cc281d5f9bf1a29d7ac08e79d7764899be8e1abc4f247875cf8db2
39b435ba73b8a740e816fa141f84d1b9d98eea1c37b59b0aeed94a205c1e424df1306b3e07b3eddbd0a94d8ae986a628acc2a93eb457d55dcebc67d799197823

$CDNENCFINISH
.ENDS COMP_0 


.SUBCKT THD_BASIC_0  VIN VOUT  
+ PARAMS: A1=1 A2=353E-6 A3=353E-6
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
dba66072656724865daad81d0b769198dc051b9a91e3562f55e03336d0061ba0ee4b01fa958f370ce4a5316a99f722437e51192624527ce4366891e1e885c871
23f81b209ce527d7197b36855ab218f42a8a2bfd4fe2703eaf193f1b96e24aebd84deecc57bef0f5616d5a9656ec2ac3fa019239cde1d81d5c249fdc134b75e9
*E_ADJUST_GAIN VOUT 0 VALUE= { V(VOUTP)*0.90909090}
$CDNENCFINISH
.ENDS THD_BASIC_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc271a8d93ed80249a
78caa60348a24a0d53ba195371f2bcb2dbe86c1f70c2d0d3d22f36355734485498459f8d9427cf6dbfb94d64dccce65cb425cc4f9b2e15f453d44eb387efa1e0
6400587cce7cd1c79b8d3130ea3e2a38f0b062208a51e23acf21098bd109a696d2e603a6aaba3a80eed94a205c1e424df1306b3e07b3eddbe3adbed052508a42
00e7e78343205e5184b1a15ace3493b904fc163d1408fe336c2f314c02bd115c29e132f0507cbf2e5442b05feec11b74ec102488afac8d9c94f258c7a007c77f
586e5476eaa3a9eac4633bb8a76cfe3e9a87dce6f28c1cabc92c652c5889c7dfaedffb309d4ac06d2c744c4029838b320afdd7f44b471c71fca3a0227cb74238
$CDNENCFINISH
.ENDS RNOISE_FREE_0 


.END

