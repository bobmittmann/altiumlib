*
*Zetex ZXMN4A06G Spice Model v3.0 Last Revised 4/12/07
*
.SUBCKT ZXMN4A06G 30 40 50
*------connections-------D-G-S
M1 6 2 5 5 Nmod L=1.16E-6 W=1.7
M2 5 2 5 6 Pmod L=1.3E-6 W=0.75
RG 4 2 1.6
RIN 2 5 1E12
RD 3 6 Rmod 0.012
RS 5 55 Rmod 0.012
RL 3 5 3E12
C1 2 5 75E-12
C2 3 4 5E-12
D1 5 3  Dbodymod
LD 3 30 1E-9
LG 4 40 2.3E-9
LS 55 50 2.3E-9
.MODEL Nmod NMOS (LEVEL=3 TOX=7.5E-8 NSUB=5E16 VTO= 1.75
+KP=1.5E-5 NFS=2E11 KAPPA=0.06 UO=650 IS=1E-15 N=10)
.MODEL Pmod PMOS (LEVEL=3 TOX=5.5E-8 NSUB=1E16
+TPG=-1 IS=1E-15 N=10)
.MODEL Dbodymod D (IS=8E-12 RS=.016 IKF=10 TRS1=1.5e-3
+CJO=250e-12  BV=44 TT=17e-9)
.MODEL Rmod RES (TC1=3.5e-3 TC2=0.8E-5)
.ENDS ZXMN4A06G
*
*$
*
*                (c)  2007 Zetex Semiconductors plc
*
*   The copyright in these models  and  the designs embodied belong
*   to Zetex Semiconductors plc (" Zetex ").  They  are  supplied
*   free of charge by Zetex for the purpose of research and design
*   and may be used or copied intact  (including this notice)  for
*   that purpose only.  All other rights are reserved. The models
*   are believed accurate but  no condition  or warranty  as to their
*   merchantability or fitness for purpose is given and no liability
*   in respect of any use is accepted by Zetex PLC, its distributors
*   or agents.
*
*   Zetex Semiconductors plc, Zetex Technology Park, Chadderton,
*   Oldham, United Kingdom, OL9 9LL