*March 21, 2005
*Doc. ID: 75256, S-50383, Rev. B
*File Name: Si3434DV_PS.txt and Si3434DV_PS.lib
.SUBCKT SI3434DV 4 1 2
M1  3 1 2 2 NMOS W=802610u L=0.50u 
M2  2 1 2 4 PMOS W=802610u L=0.50u
R1  4 3     RTEMP 14E-3
CGS 1 2     380E-12
DBD 2 4     DBD
**************************************************************************
.MODEL  NMOS       NMOS (  LEVEL  = 3               TOX    = 3E-8
+ RS     = 6.5E-3          RD     = 0               NSUB   = 1.85E17   
+ kp     = 3.1E-5          UO     = 650             
+ VMAX   = 0               XJ     = 5E-7            KAPPA  = 2E-2
+ ETA    = 1E-4            TPG    = 1  
+ IS     = 0               LD     = 0                             
+ CGSO   = 0               CGDO   = 0               CGBO   = 0 
+ NFS    = 0.8E12          DELTA  = 0.1)
*************************************************************************
.MODEL  PMOS       PMOS (LEVEL    = 3               TOX    = 3E-8
+NSUB    = 5E16            TPG    = -1)           
*************************************************************************
.MODEL DBD D (CJO=270E-12  VJ=.38   M=0.3
+RS=0.1 FC=0.1 IS=1E-12 TT=4E-8 N=1 BV=30.5)
*************************************************************************
.MODEL RTEMP RES (TC1=6E-3   TC2=5.5E-6)
*************************************************************************
.ENDS
 
