* OPA365 SPICE MACROMODEL
*          
*   Rev. A    4 August 2006, by W.K. SANDS
*
*   Rev. B    4 August 2006, by NEIL ALBAUGH: ADDED HEADER TEXT & EDITED TEXT
*
*
*     This macromodel has been optimized to model the AC, DC, and transient response performance within 
*     the device data sheet specified limits. 
*     Correct operation of this macromodel has been verified on MicroSim P-Spice ver. 8.0, DesignSoft TINA, and on 
*     PENZAR Development TopSPICE ver. 6.82d. For help with other analog simulation software, 
*     please consult your software supplier. 
*
*  
*   Copyright 2006 by Texas Instruments Corporation
*
* MODEL TEMPERATURE RANGE IS -40 C TO +125 C, NOT ALL PARAMETERS ACCURATELY TRACK THOSE OF AN ACTUAL OPA365 
* OVER THE FULL TEMPERATURE RANGE BUT ARE AS CLOSE AS PRACTICAL
*
* END NOTES
*
* BEGIN MODEL OPA365
*
* BEGIN MODEL FEATURES
*
* OPEN LOOP GAIN AND PHASE
* INPUT VOLTAGE NOISE
* INPUT CURRENT NOISE
* INPUT BIAS CURRENT
* INPUT CAPACITANCE
* INPUT COMMON MODE VOLTAGE RANGE
* INPUT CLAMPS TO RAILS
* CMRR WITH FREQUENCY EFFECTS
* PSRR WITH FREQUENCY EFFECTS
* SLEW RATE
* SETTLING TIME
* OVERLOAD RECOVERY TIME
* QUIESCENT CURRENT
* QUIESCENT CURRENT VS VOLTAGE
* RAIL TO RAIL OUTPUT STAGE
* HIGH CLOAD EFFECTS
* CLASS AB BIAS IN OUTPUT STAGE
* OUTPUT CURRENT THROUGH SUPPLIES
* OUTPUT CURRENT LIMITING
* OUTPUT CLAMPS TO RAILS
* OUTPUT SWING VS OUTPUT CURRENT
*
* END MODEL FEATURES
*
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   4   5  2  1
*
.SUBCKT OPA365 3 4 5 2 1
*
Q23 6 7 8 QNL
R211 9 10 2
R212 11 10 2
R213 7 12 1E3
R214 13 14 1E3
R215 15 5 8
R216 2 16 8
R218 17 18 250
R219 19 20 8
R220 8 21 8
D33 22 5 DD
D34 2 22 DD
D35 23 0 DIN
D36 24 0 DIN
I29 0 23 0.1E-3
I30 0 24 0.1E-3
E72 8 0 2 0 1
E73 20 0 5 0 1
D37 25 0 DVN
D38 26 0 DVN
I31 0 25 0.1E-3
I32 0 26 0.1E-3
E74 27 4 25 26 0.32
G25 28 4 23 24 1.75E-6
R221 2 5 5E3
E75 29 0 20 0 1
E76 30 0 8 0 1
E77 31 0 32 0 1
R223 29 33 1E5
R224 30 34 1E5
R225 31 35 1E5
R226 0 33 10
R227 0 34 10
R228 0 35 10
E78 36 3 35 0 0.003
R229 37 32 1E3
R230 32 38 1E3
C50 29 33 1E-12
C51 30 34 1E-12
C52 31 35 5E-9
E79 39 36 34 0 -0.15
E80 28 39 33 0 0.15
E81 40 8 20 8 0.5
D39 17 20 DD
D40 8 17 DD
M61 41 42 16 16 NOUT L=3U W=1600U
M62 43 44 15 15 POUT L=3U W=1600U
M63 45 45 19 19 POUT L=3U W=1600U
M64 46 47 9 9 PIN L=3U W=440U
M65 48 49 11 11 PIN L=3U W=440U
M66 50 50 21 21 NOUT L=3U W=1600U
R231 51 44 100
R232 52 42 100
G26 17 40 53 40 0.2E-3
R233 40 17 20E6
C53 18 22 4.2E-12
R234 8 46 3E3
R235 8 48 3E3
C54 46 48 0.08E-12
C55 28 0 6E-12
C56 27 0 6E-12
C57 22 0 5E-12
D41 42 6 DD
D42 54 44 DD
Q24 54 14 20 QPL
V93 28 55 75E-6
M67 56 57 20 20 PIN L=6U W=500U
E82 38 0 28 0 1
E83 37 0 4 0 1
M68 57 57 20 20 PIN L=6U W=500U
V95 56 10 -0.9
R236 22 43 8
R237 41 22 8
J9 20 28 20 JI
J10 20 27 20 JI
J11 27 58 27 JI
J12 28 58 28 JI
C58 28 27 0.35E-12
E84 59 40 48 46 1
R238 59 53 1E4
C59 53 40 0.08E-12
G27 60 40 17 40 -1E-3
G28 40 61 17 40 1E-3
G29 40 62 50 8 1E-3
G30 63 40 20 45 1E-3
D43 63 60 DD
D44 61 62 DD
R239 60 63 100E6
R240 62 61 100E6
R241 63 20 1E3
R242 8 62 1E3
E85 20 51 20 63 1
E86 52 8 62 8 1
R243 61 40 1E6
R244 62 40 1E6
R245 40 63 1E6
R246 40 60 1E6
R247 0 64 1E6
R248 39 28 1E9
R249 36 39 1E9
R250 3 36 1E9
R251 4 27 1E9
R252 40 53 1E9
R253 51 20 1E9
R254 8 52 1E9
R255 32 0 1E9
G32 57 8 64 0 181E-6
G33 45 50 64 0 490E-6
I35 5 2 3.15E-3
L5 22 1 0.4E-9
R265 22 1 400
R269 45 20 1E8
R270 8 50 1E8
R271 15 44 1E8
R272 42 22 1E8
G36 27 0 65 0 23E-12
I42 27 0 200E-15
I47 0 66 1M
D46 66 0 DD
V113 66 67 0.655
R311 0 67 1E6
E94 68 0 67 0 -571
R312 0 68 1E6
G37 28 0 65 0 23E-12
I49 28 0 200E-15
V119 69 68 -73
D47 69 65 DD
R313 0 65 1E6
R315 47 55 100
R316 27 49 100
V120 58 8 0.3
R317 57 20 1E9
V121 64 0 1
R380 17 22 1E9
E115 12 8 16 8 1.5
E116 20 13 5 15 1.5
.MODEL DVN D KF=8E-14 IS=1E-16
.MODEL DIN D
.MODEL DD D
.MODEL JI NJF IS=1E-18
.MODEL QPL PNP
.MODEL QNL NPN
.MODEL POUT PMOS KP=200U VTO=-0.7
.MODEL NOUT NMOS KP=200U VTO=0.7
.MODEL PIN PMOS KP=200U VTO=-0.7
.ENDS
* END MODEL OPA365
