.SUBCKT BCM62B 1 2 3 4

*
* Pin 1: Collector;Base  TR2; TR1 and TR2
* Pin 2: Collector       TR1
* Pin 3: Emitter         TR1
* Pin 4: Emitter         TR2
*

*  C B E 
Q1 2 1 3 QBCM62B
*  C B E 
Q2 1 1 4 QBCM62B

*
**********************************************************
*
* BCM62B
*
* NXP Semiconductors
*
* Matched double PNP/PNP transistor
* IC   = 100 mA
* VCEO = 45 V 
* hFE  = 200 - 450 @ 5V/2mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 143
* 
* Package Pin 1:   Collector;Base   	TR2; TR1 and TR2
* Package Pin 2:   Collector        	TR1
* Package Pin 3;4: Emitter          	TR1;TR2
*
*
* Extraction date (week/year): 14/2006
* Simulator: Spice 2        
*
**********************************************************
*#
* Please note: The following model is to be used twice in 
* schematic due to equality of both transistors.
*
.MODEL QBCM62B PNP
+     IS = 2.014E-14 
+     NF = 0.9974 
+     ISE = 6.578E-15 
+     NE = 1.45 
+     BF = 315.3 
+     IKF = 0.079 
+     VAF = 39.15 
+     NR = 0.9952 
+     ISC = 1.633E-14 
+     NC = 1.15 
+     BR = 8.68 
+     IKR = 0.09 
+     VAR = 9.5 
+     RB = 10 
+     IRB = 5E-06 
+     RBM = 5E-06 
+     RE = 0.663 
+     RC = 0.718 
+     XTB = 0 
+     EG = 1.11 
+     XTI = 3 
+     CJE = 1.135E-11 
+     VJE = 0.7071 
+     MJE = 0.3808 
+     TF = 6.546E-10 
+     XTF = 5.387 
+     VTF = 6.245 
+     ITF = 0.2108 
+     PTF = 0 
+     CJC = 6.395E-12 
+     VJC = 0.4951 
+     MJC = 0.44 
+     XCJC = 0.6288 
+     TR = 5.5E-08 
+     CJS = 0 
+     VJS = 0.75 
+     MJS = 0.333  
+     FC = 0.9059
*##
*

.ENDS

