*TITLE=ZXCT1010 MACROMODEL
*ORIGIN=DZSL_AG_GS
*SIMULATOR=DIODES, SIMETRIX and PSPICE
*DATE=14th July 2010
*VERSION=1
*PIN_ORDER     2:GND, 3:OUT, 4:S+, 5:S-   (Pin 1 is NC)
*
.subckt ZXCT1010 GND OUT S+ S-
* pins------------2---3--4--5
*
R1  S- FILT  100k      ;input filter
C1  S+ FILT  20p       ;input filter
R2  S+ GND  1Meg       ;quiescent current at 5V
*  Output as a voltage: first part of expression limits resonse to zero for negative input
*  tanh function limits output when supply is less than 1.1V above Vout
E1  E1OUT GND VALUE={ max(V(S+)-V(FILT),0)*tanh( 20*max(V(S-)-1.1-V(OUT),0) ) }
R3  E1OUT GND 1Meg
*  Transconductance = 1/100 A/V, with temperature dependence
G1  S+  OUT VALUE={(V(E1OUT) - V(GND))*(1/100)*(1.01-0.0003*TEMP-6e-6*(TEMP**2)-5e-8*(TEMP**3)+2.7e-10*(TEMP**4))}
.ends ZXCT1010
*
*
*                (c)  2010 Diodes Inc
*
*   The copyright in these models  and  the designs embodied belong
*   to Diodes Incorporated (" Zetex ").  They  are  supplied
*   free of charge by Zetex for the purpose of research and design
*   and may be used or copied intact  (including this notice)  for
*   that purpose only.  All other rights are reserved.  The models
*   are believed accurate but no condition  or warranty  as to their
*   merchantability or fitness for purpose is given and no liability
*   in respect of any use is accepted by Diodes Incorporated, its distributors
*   or agents.
*
*   Diodes Zetex Semiconductors Ltd, Zetex Technology Park, Chadderton,
*   Oldham, United Kingdom, OL9 9LL
*
*
